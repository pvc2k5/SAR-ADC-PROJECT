** sch_path: /home/tien/gf180ex/ADC_SAR.sch
**.subckt ADC_SAR Valid VOCP VOCN Vinp Vinn VDD Vinp S1 Vpositive Vnegative Vcm Vrefp Vrefn Vrefn Vrefp Vcm Vrefp Vcm Vrefn S0 E
*+ Vinn S1 S0 E VDD VDD VDD S1 S0 E
*.opin Valid
*.opin VOCP
*.opin VOCN
*.ipin Vinp
*.ipin Vinn
*.iopin VDD
*.ipin Vinp
*.ipin S1
*.opin Vpositive
*.opin Vnegative
*.ipin Vcm
*.ipin Vrefp
*.ipin Vrefn
*.ipin Vrefn
*.ipin Vrefp
*.ipin Vcm
*.ipin Vrefp
*.ipin Vcm
*.ipin Vrefn
*.ipin S0
*.ipin E
*.ipin Vinn
*.ipin S1
*.ipin S0
*.ipin E
*.iopin VDD
*.iopin VDD
*.iopin VDD
*.ipin S1
*.ipin S0
*.ipin E
x1 VDD VOCP Vpositive Vnegative Valid VOCN nCLK CLK GND cp2
XC63 Vpositive net8 cap_mim_1f0fF c_width=1.182e-6 c_length=2.644e-6 m=1
XC126 Vnegative net19 cap_mim_1f0fF c_width=1.182e-6 c_length=2.644e-6 m=1
x4 net2 Vpositive 16C
x5 Vpositive net1 8C
x6 net23 Vpositive 4C
x7 net22 Vpositive 2C
x8 net21 Vpositive C
x9 net7 net8 16C
x10 net8 net6 8C
x11 net5 net8 4C
x12 net4 net8 2C
x13 net3 net8 C
x14 net13 Vnegative 16C
x15 Vnegative net12 8C
x16 net11 Vnegative 4C
x17 net10 Vnegative 2C
x18 net9 Vnegative C
x19 net18 net19 16C
x20 net19 net17 8C
x21 net16 net19 4C
x22 net15 net19 2C
x23 net14 net19 C
V11 VDD GND 3.3
V12 CLK GND PULSE(0 3.3 0 0.5n 0.5n 40n 100n)

V13 nCLK GND PULSE(3.3 0 0 0.5n 0.5n 40n 100n)

V4 Vinp net20 SIN(0.9 0.9 10Meg) DC 0
V5 net20 GND 0
V1 Vinn GND 1.5
x24 VDD Vinp E CLK nCLK Vcm net2 Vrefp Vrefn S0 S1 GND MUX4_1
x2 VDD Vinp E CLK nCLK Vcm net1 Vrefp Vrefn S0 S1 GND MUX4_1
x25 VDD Vinp CLK CLK nCLK Vcm net23 Vrefp Vrefn S0 S1 GND MUX4_1
x26 VDD Vinp E CLK nCLK Vcm net22 Vrefp Vrefn S0 S1 GND MUX4_1
x27 VDD Vinp E CLK nCLK Vcm net21 Vrefp Vrefn S0 S1 GND MUX4_1
x28 VDD Vinp E CLK nCLK Vcm net7 Vrefp Vrefn S0 S1 GND MUX4_1
x29 VDD Vinp E CLK nCLK Vcm net6 Vrefp Vrefn S0 S1 GND MUX4_1
x30 VDD Vinp E CLK nCLK Vcm net5 Vrefp Vrefn S0 S1 GND MUX4_1
x31 VDD Vinp E CLK nCLK Vcm net4 Vrefp Vrefn S0 S1 GND MUX4_1
x32 VDD Vinp E CLK nCLK Vcm net3 Vrefp Vrefn S0 S1 GND MUX4_1
x3 VDD Vinn E CLK nCLK Vcm net13 Vrefp Vrefn S0 S1 GND MUX4_1N
x33 VDD Vinn E CLK nCLK Vcm net12 Vrefp Vrefn S0 S1 GND MUX4_1N
x34 VDD Vinn E CLK nCLK Vcm net11 Vrefp Vrefn S0 S1 GND MUX4_1N
x35 VDD Vinn E CLK nCLK Vcm net10 Vrefp Vrefn S0 S1 GND MUX4_1N
x36 VDD Vinn E CLK nCLK Vcm net9 Vrefp Vrefn S0 S1 GND MUX4_1N
x37 VDD Vinn E CLK nCLK Vcm net18 Vrefp Vrefn S0 S1 GND MUX4_1N
x38 VDD Vinn E CLK nCLK Vcm net17 Vrefp Vrefn S0 S1 GND MUX4_1N
x39 VDD Vinn E CLK nCLK Vcm net16 Vrefp Vrefn S0 S1 GND MUX4_1N
x40 VDD Vinn E CLK nCLK Vcm net15 Vrefp Vrefn S0 S1 GND MUX4_1N
x41 VDD Vinn E CLK nCLK Vcm net14 Vrefp Vrefn S0 S1 GND MUX4_1N
V2 Vrefp GND 3.3
V3 Vcm GND 1.65
V6 Vrefn GND 0
V7 S0 GND PULSE(0 3.3 0 0.5n 0.5n 40n 100n)


V8 S1 GND PULSE(0 3.3 0 0.5n 0.5n 100n 200n)

V9 E GND 3.3
**** begin user architecture code

.tran 0.01n 1u
.temp 25
.save all



.include /home/tien/conda-gf180mcu-env/envs/gf180mcu-env/share/pdk/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/tien/conda-gf180mcu-env/envs/gf180mcu-env/share/pdk/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical
.lib /home/tien/conda-gf180mcu-env/envs/gf180mcu-env/share/pdk/gf180mcuC/libs.tech/ngspice/smbb000149.ngspice typical
.lib /home/tien/conda-gf180mcu-env/envs/gf180mcu-env/share/pdk/gf180mcuC/libs.tech/ngspice/sm141064.ngspice cap_mim
.lib /home/tien/conda-gf180mcu-env/envs/gf180mcu-env/share/pdk/gf180mcuC/libs.tech/ngspice/sm141064.ngspice mimcap_typical
.lib /home/tien/conda-gf180mcu-env/envs/gf180mcu-env/share/pdk/gf180mcuC/libs.tech/ngspice/sm141064.ngspice res_typical
.lib /home/tien/conda-gf180mcu-env/envs/gf180mcu-env/share/pdk/gf180mcuC/libs.tech/ngspice/sm141064.ngspice moscap_typical

**** end user architecture code
**.ends

* expanding   symbol:  cp2.sym # of pins=9
** sym_path: /home/tien/gf180ex/cp2.sym
** sch_path: /home/tien/gf180ex/cp2.sch
.subckt cp2 VP VOCP VDP VDN Valid VOCN nCLK CLK VN
*.iopin VP
*.iopin CLK
*.iopin nCLK
*.ipin VDP
*.ipin VDN
*.opin Valid
*.opin VOCP
*.opin VOCN
*.iopin VN
XM1 net4 CLK VP VP pfet_03v3 L=0.28u W=3.9u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM2 net3 CLK VP VP pfet_03v3 L=0.28u W=3.9u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM3 net2 net7 VP VP pfet_03v3 L=0.28u W=16u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM4 net1 net6 VP VP pfet_03v3 L=0.28u W=16u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM5 net7 net4 net1 VP pfet_03v3 L=0.28u W=16u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM6 net6 net3 net2 VP pfet_03v3 L=0.28u W=16u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM7 net3 VDP net5 GND nfet_03v3 L=0.28u W=0.9u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM8 net4 VDN net5 GND nfet_03v3 L=0.28u W=0.9u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM9 net5 CLK VN VN nfet_03v3 L=0.28u W=10u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM10 net7 nCLK VN VN nfet_03v3 L=0.28u W=3.1u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM11 net7 net6 VN VN nfet_03v3 L=0.28u W=6.2u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM12 net6 net7 VN VN nfet_03v3 L=0.28u W=6.2u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM13 net6 nCLK VN VN nfet_03v3 L=0.28u W=3.1u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
x3 VP Valid VOCP VOCN VN NAND
x1 VP VOCP net6 VN inverter
x2 VP VOCN net7 VN inverter
.ends


* expanding   symbol:  16C.sym # of pins=2
** sym_path: /home/tien/gf180ex/16C.sym
** sch_path: /home/tien/gf180ex/16C.sch
.subckt 16C bottom_plate top_plate
*.iopin bottom_plate
*.iopin top_plate
XC1 bottom_plate top_plate cap_mim_1f0fF c_width=1.182e-6 c_length=2.644e-6 m=1
XC2 bottom_plate top_plate cap_mim_1f0fF c_width=1.182e-6 c_length=2.644e-6 m=1
XC3 bottom_plate top_plate cap_mim_1f0fF c_width=1.182e-6 c_length=2.644e-6 m=1
XC4 bottom_plate top_plate cap_mim_1f0fF c_width=1.182e-6 c_length=2.644e-6 m=1
XC5 bottom_plate top_plate cap_mim_1f0fF c_width=1.182e-6 c_length=2.644e-6 m=1
XC6 bottom_plate top_plate cap_mim_1f0fF c_width=1.182e-6 c_length=2.644e-6 m=1
XC7 bottom_plate top_plate cap_mim_1f0fF c_width=1.182e-6 c_length=2.644e-6 m=1
XC8 bottom_plate top_plate cap_mim_1f0fF c_width=1.182e-6 c_length=2.644e-6 m=1
XC9 bottom_plate top_plate cap_mim_1f0fF c_width=1.182e-6 c_length=2.644e-6 m=1
XC10 bottom_plate top_plate cap_mim_1f0fF c_width=1.182e-6 c_length=2.644e-6 m=1
XC11 bottom_plate top_plate cap_mim_1f0fF c_width=1.182e-6 c_length=2.644e-6 m=1
XC12 bottom_plate top_plate cap_mim_1f0fF c_width=1.182e-6 c_length=2.644e-6 m=1
XC13 bottom_plate top_plate cap_mim_1f0fF c_width=1.182e-6 c_length=2.644e-6 m=1
XC14 bottom_plate top_plate cap_mim_1f0fF c_width=1.182e-6 c_length=2.644e-6 m=1
XC15 bottom_plate top_plate cap_mim_1f0fF c_width=1.182e-6 c_length=2.644e-6 m=1
XC16 bottom_plate top_plate cap_mim_1f0fF c_width=1.182e-6 c_length=2.644e-6 m=1
.ends


* expanding   symbol:  8C.sym # of pins=2
** sym_path: /home/tien/gf180ex/8C.sym
** sch_path: /home/tien/gf180ex/8C.sch
.subckt 8C top_plate bottom_plate
*.iopin bottom_plate
*.iopin top_plate
XC2 bottom_plate top_plate cap_mim_1f0fF c_width=1.182e-6 c_length=2.644e-6 m=1
XC3 bottom_plate top_plate cap_mim_1f0fF c_width=1.182e-6 c_length=2.644e-6 m=1
XC4 bottom_plate top_plate cap_mim_1f0fF c_width=1.182e-6 c_length=2.644e-6 m=1
XC5 bottom_plate top_plate cap_mim_1f0fF c_width=1.182e-6 c_length=2.644e-6 m=1
XC6 bottom_plate top_plate cap_mim_1f0fF c_width=1.182e-6 c_length=2.644e-6 m=1
XC7 bottom_plate top_plate cap_mim_1f0fF c_width=1.182e-6 c_length=2.644e-6 m=1
XC8 bottom_plate top_plate cap_mim_1f0fF c_width=1.182e-6 c_length=2.644e-6 m=1
XC1 bottom_plate top_plate cap_mim_1f0fF c_width=1.182e-6 c_length=2.644e-6 m=1
.ends


* expanding   symbol:  4C.sym # of pins=2
** sym_path: /home/tien/gf180ex/4C.sym
** sch_path: /home/tien/gf180ex/4C.sch
.subckt 4C bottom_plate top_plate
*.iopin top_plate
*.iopin bottom_plate
XC5 bottom_plate top_plate cap_mim_1f0fF c_width=1.182e-6 c_length=2.644e-6 m=1
XC6 bottom_plate top_plate cap_mim_1f0fF c_width=1.182e-6 c_length=2.644e-6 m=1
XC7 bottom_plate top_plate cap_mim_1f0fF c_width=1.182e-6 c_length=2.644e-6 m=1
XC8 bottom_plate top_plate cap_mim_1f0fF c_width=1.182e-6 c_length=2.644e-6 m=1
.ends


* expanding   symbol:  2C.sym # of pins=2
** sym_path: /home/tien/gf180ex/2C.sym
** sch_path: /home/tien/gf180ex/2C.sch
.subckt 2C bottom_plate top_plate
*.iopin top_plate
*.iopin bottom_plate
XC5 bottom_plate top_plate cap_mim_1f0fF c_width=1.182e-6 c_length=2.644e-6 m=1
XC6 bottom_plate top_plate cap_mim_1f0fF c_width=1.182e-6 c_length=2.644e-6 m=1
.ends


* expanding   symbol:  C.sym # of pins=2
** sym_path: /home/tien/gf180ex/C.sym
** sch_path: /home/tien/gf180ex/C.sch
.subckt C bottom_plate top_plate
*.iopin bottom_plate
*.iopin top_plate
XC5 bottom_plate top_plate cap_mim_1f0fF c_width=1.182e-6 c_length=2.644e-6 m=1
.ends


* expanding   symbol:  MUX4_1.sym # of pins=12
** sym_path: /home/tien/gf180ex/MUX4_1.sym
** sch_path: /home/tien/gf180ex/MUX4_1.sch
.subckt MUX4_1 VP Vinp E CLK nCLK Vcm Vout Vrefp Vrefn S0 S1 VN
*.iopin VP
*.ipin E
*.opin Vout
*.ipin Vcm
*.ipin Vrefp
*.ipin Vrefn
*.ipin S0
*.ipin S1
*.ipin Vinp
*.ipin CLK
*.ipin nCLK
*.iopin VN
x1 VP net2 E net1 net6 net7 VN And
x2 VP net3 E Vcm net6 net8 VN And
x3 VP net4 E Vrefp net9 net7 VN And
x4 VP net5 E Vrefn net9 net8 VN And
x5 VP CLK net1 nCLK Vinp VN sample2
x6 VP net2 net3 net4 net5 Vout VN OR
x7 VP net6 S0 VN inverter
x8 VP net9 net6 VN inverter
x9 VP net7 S1 VN inverter
x10 VP net8 net7 VN inverter
.ends


* expanding   symbol:  MUX4_1N.sym # of pins=12
** sym_path: /home/tien/gf180ex/MUX4_1N.sym
** sch_path: /home/tien/gf180ex/MUX4_1N.sch
.subckt MUX4_1N VP Vinn E CLK nCLK Vcm Vout Vrefp Vrefn S0 S1 VN
*.iopin VP
*.ipin E
*.opin Vout
*.ipin Vcm
*.ipin Vrefp
*.ipin Vrefn
*.ipin S0
*.ipin S1
*.ipin Vinn
*.ipin CLK
*.ipin nCLK
*.iopin VN
x1 VP net2 E net1 net6 net7 VN And
x2 VP net3 E Vcm net6 net8 VN And
x3 VP net4 E Vrefp net9 net7 VN And
x4 VP net5 E Vrefn net9 net8 VN And
x6 VP net2 net3 net4 net5 Vout VN OR
x7 VP net6 S0 VN inverter
x8 VP net9 net6 VN inverter
x9 VP net7 S1 VN inverter
x10 VP net8 net7 VN inverter
x11 VP CLK net1 nCLK Vinn VN sa2_n
.ends


* expanding   symbol:  NAND.sym # of pins=5
** sym_path: /home/tien/gf180ex/NAND.sym
** sch_path: /home/tien/gf180ex/NAND.sch
.subckt NAND VP Vout A B VN
*.iopin VP
*.ipin A
*.ipin B
*.opin Vout
*.iopin VN
XM1 Vout B VP VP pfet_03v3 L=0.28u W=2.8u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM2 Vout A VP VP pfet_03v3 L=0.28u W=2.8u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM3 Vout A net1 VN nfet_03v3 L=0.28u W=1u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM4 net1 B VN VN nfet_03v3 L=0.28u W=1u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  inverter.sym # of pins=4
** sym_path: /home/tien/gf180ex/inverter.sym
** sch_path: /home/tien/gf180ex/inverter.sch
.subckt inverter Vp Vout Vin VN
*.iopin Vp
*.ipin Vin
*.opin Vout
*.iopin VN
XM1 Vout Vin Vp Vp pfet_03v3 L=0.28u W=2.8u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM2 Vout Vin VN VN nfet_03v3 L=0.28u W=1u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  And.sym # of pins=7
** sym_path: /home/tien/gf180ex/And.sym
** sch_path: /home/tien/gf180ex/And.sch
.subckt And VP Vout A B C D VN
*.ipin A
*.ipin B
*.ipin C
*.ipin D
*.iopin VP
*.iopin VN
*.opin Vout
XM1 net1 A net3 VN nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM2 net3 B net4 VN nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM3 net4 C net5 VN nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM4 net5 D VN VN nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM5 net2 D VP VP pfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM6 net2 C VP VP pfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM7 net2 B VP VP pfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM8 net1 A VP VP pfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
x1 VP Vout net2 VN inverter
.ends


* expanding   symbol:  sample2.sym # of pins=6
** sym_path: /home/tien/gf180ex/sample2.sym
** sch_path: /home/tien/gf180ex/sample2.sch
.subckt sample2 VP CLK Vout nCLK Vinp VN
*.ipin Vinp
*.opin Vout
*.iopin VP
*.iopin CLK
*.iopin nCLK
*.iopin VN
XM1 net4 CLK VP VP pfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM2 VP net2 net1 net1 pfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM3 net2 net4 net1 net1 pfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM4 net2 VP net3 VN nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM5 net3 nCLK VN VN nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM6 net4 CLK net5 VN nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM7 net4 net2 net5 VN nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM8 Vinp net2 net5 VN nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM9 Vout net2 Vinp VN nfet_03v3 L=0.28u W=0.39u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XC1 net1 net5 cap_mim_1f0fF c_width=100e-6 c_length=10e-6 m=1
XC2 Vout VN cap_mim_1f0fF c_width=3e-6 c_length=1e-6 m=1
XM10 net5 nCLK VN VN nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  OR.sym # of pins=7
** sym_path: /home/tien/gf180ex/OR.sym
** sch_path: /home/tien/gf180ex/OR.sch
.subckt OR VP A B C D Vout VN
*.ipin A
*.ipin B
*.ipin C
*.ipin D
*.opin Vout
*.iopin VP
*.iopin VN
XM1 net2 A VN VN nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM2 net2 B VN VN nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM3 net2 C VN VN nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM4 net1 D VN VN nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM5 net1 D net3 VP pfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM6 net3 C net4 VP pfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM7 net4 B net5 VP pfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM8 net5 A VP VP pfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
x1 VP Vout net2 VN inverter
.ends


* expanding   symbol:  sa2_n.sym # of pins=6
** sym_path: /home/tien/gf180ex/sa2_n.sym
** sch_path: /home/tien/gf180ex/sa2_n.sch
.subckt sa2_n VP CLK Vout nCLK Vinn VN
*.ipin Vinn
*.opin Vout
*.iopin VP
*.iopin CLK
*.iopin nCLK
*.iopin VN
XM1 net4 CLK VP VP pfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM2 VP net2 net1 net1 pfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM3 net2 net4 net1 net1 pfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM4 net2 VP net3 VN nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM5 net3 nCLK VN VN nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM6 net4 CLK net5 VN nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM7 net4 net2 net5 VN nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM8 Vinn net2 net5 VN nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM9 Vout net2 Vinn VN nfet_03v3 L=0.28u W=0.39u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XC1 net1 net5 cap_mim_1f0fF c_width=100e-6 c_length=10e-6 m=1
XC2 Vout VN cap_mim_1f0fF c_width=3e-6 c_length=1e-6 m=1
XM10 net5 nCLK VN VN nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
.ends

.GLOBAL GND
.end
