module adc_core_digital (a_clk_dig_in,
    a_comparator_in,
    a_conv_finished_osr_out,
    a_enable_loop_out,
    a_nmatrix_c0_out_n,
    a_pmatrix_c0_out_n,
    a_rst_n,
    a_sample_matrix_out,
    a_sample_matrix_out_n,
    a_sample_switch_out,
    a_sample_switch_out_n,
    a_config_1_in,
    a_config_2_in,
    a_nmatrix_bincap_out_n,
    a_nmatrix_col_out,
    a_nmatrix_col_out_n,
    a_nmatrix_row_out_n,
    a_nmatrix_rowoff_out_n,
    a_nmatrix_rowon_out_n,
    a_pmatrix_bincap_out_n,
    a_pmatrix_col_out,
    a_pmatrix_col_out_n,
    a_pmatrix_row_out_n,
    a_pmatrix_rowoff_out_n,
    a_pmatrix_rowon_out_n,
    a_result_out);
 input a_clk_dig_in;
 input a_comparator_in;
 output a_conv_finished_osr_out;
 output a_enable_loop_out;
 output a_nmatrix_c0_out_n;
 output a_pmatrix_c0_out_n;
 input a_rst_n;
 output a_sample_matrix_out;
 output a_sample_matrix_out_n;
 output a_sample_switch_out;
 output a_sample_switch_out_n;
 input [9:0] a_config_1_in;
 input [9:0] a_config_2_in;
 output [2:0] a_nmatrix_bincap_out_n;
 output [12:0] a_nmatrix_col_out;
 output [12:0] a_nmatrix_col_out_n;
 output [9:0] a_nmatrix_row_out_n;
 output [9:0] a_nmatrix_rowoff_out_n;
 output [9:0] a_nmatrix_rowon_out_n;
 output [2:0] a_pmatrix_bincap_out_n;
 output [12:0] a_pmatrix_col_out;
 output [12:0] a_pmatrix_col_out_n;
 output [9:0] a_pmatrix_row_out_n;
 output [9:0] a_pmatrix_rowoff_out_n;
 output [9:0] a_pmatrix_rowon_out_n;
 output [9:0] a_result_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0373_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0383_;
 wire _0384_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire net10;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire net9;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire net8;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire net7;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire clknet_2_0__leaf_a_clk_dig_in;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire clknet_0_a_clk_dig_in;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire clknet_2_3__leaf_a_clk_dig_in;
 wire clknet_2_1__leaf_a_clk_dig_in;
 wire clknet_2_2__leaf_a_clk_dig_in;
 wire \cnb.average_counter_r[0] ;
 wire \cnb.average_counter_r[1] ;
 wire \cnb.average_counter_r[2] ;
 wire \cnb.average_counter_r[3] ;
 wire \cnb.average_counter_r[4] ;
 wire \cnb.average_sum_r[0] ;
 wire \cnb.average_sum_r[1] ;
 wire \cnb.average_sum_r[2] ;
 wire \cnb.average_sum_r[3] ;
 wire \cnb.average_sum_r[4] ;
 wire \cnb.conv_finished_r ;
 wire net6;
 wire net5;
 wire net4;
 wire \cnb.data_register_r[3] ;
 wire \cnb.data_register_r[4] ;
 wire \cnb.data_register_r[5] ;
 wire \cnb.data_register_r[6] ;
 wire \cnb.data_register_r[7] ;
 wire \cnb.data_register_r[8] ;
 wire \cnb.data_register_r[9] ;
 wire \cnb.is_holding_result_w ;
 wire \cnb.next_average_counter_w[0] ;
 wire \cnb.next_average_counter_w[1] ;
 wire \cnb.next_average_counter_w[2] ;
 wire \cnb.next_average_counter_w[3] ;
 wire \cnb.next_average_counter_w[4] ;
 wire \cnb.next_average_sum_w[0] ;
 wire \cnb.next_average_sum_w[1] ;
 wire \cnb.next_average_sum_w[2] ;
 wire \cnb.next_average_sum_w[3] ;
 wire \cnb.next_average_sum_w[4] ;
 wire \cnb.result_out[0] ;
 wire \cnb.result_out[1] ;
 wire \cnb.result_out[2] ;
 wire \cnb.result_out[3] ;
 wire \cnb.result_out[4] ;
 wire \cnb.result_out[5] ;
 wire \cnb.result_out[6] ;
 wire \cnb.result_out[7] ;
 wire \cnb.result_out[8] ;
 wire \cnb.result_out[9] ;
 wire \cnb.result_strobe_w ;
 wire \cnb.sampled_avg_control_r[0] ;
 wire \cnb.sampled_avg_control_r[1] ;
 wire \cnb.sampled_avg_control_r[2] ;
 wire \cnb.shift_register_r[10] ;
 wire \cnb.shift_register_r[11] ;
 wire \cnb.shift_register_r[12] ;
 wire \cnb.shift_register_r[13] ;
 wire \cnb.shift_register_r[14] ;
 wire \cnb.shift_register_r[2] ;
 wire \cnb.shift_register_r[3] ;
 wire \cnb.shift_register_r[4] ;
 wire \cnb.shift_register_r[5] ;
 wire \cnb.shift_register_r[6] ;
 wire \cnb.shift_register_r[7] ;
 wire \cnb.shift_register_r[8] ;
 wire \cnb.shift_register_r[9] ;
 wire \osr.data_valid_r ;
 wire \osr.is_last_sample ;
 wire \osr.next_result_w[0] ;
 wire \osr.next_result_w[10] ;
 wire \osr.next_result_w[11] ;
 wire \osr.next_result_w[12] ;
 wire \osr.next_result_w[13] ;
 wire \osr.next_result_w[14] ;
 wire \osr.next_result_w[15] ;
 wire \osr.next_result_w[1] ;
 wire \osr.next_result_w[2] ;
 wire \osr.next_result_w[3] ;
 wire \osr.next_result_w[4] ;
 wire \osr.next_result_w[5] ;
 wire \osr.next_result_w[6] ;
 wire \osr.next_result_w[7] ;
 wire \osr.next_result_w[8] ;
 wire \osr.next_result_w[9] ;
 wire \osr.next_sample_count_w[0] ;
 wire \osr.next_sample_count_w[1] ;
 wire \osr.next_sample_count_w[2] ;
 wire \osr.next_sample_count_w[3] ;
 wire \osr.next_sample_count_w[4] ;
 wire \osr.next_sample_count_w[5] ;
 wire \osr.next_sample_count_w[6] ;
 wire \osr.next_sample_count_w[7] ;
 wire \osr.next_sample_count_w[8] ;
 wire \osr.osr_mode_r[0] ;
 wire \osr.osr_mode_r[1] ;
 wire \osr.osr_mode_r[2] ;
 wire \osr.result_r[0] ;
 wire \osr.result_r[10] ;
 wire \osr.result_r[11] ;
 wire \osr.result_r[12] ;
 wire \osr.result_r[13] ;
 wire \osr.result_r[14] ;
 wire \osr.result_r[15] ;
 wire \osr.result_r[1] ;
 wire \osr.result_r[2] ;
 wire \osr.result_r[3] ;
 wire \osr.result_r[4] ;
 wire \osr.result_r[5] ;
 wire \osr.result_r[6] ;
 wire \osr.result_r[7] ;
 wire \osr.result_r[8] ;
 wire \osr.result_r[9] ;
 wire \osr.sample_count_r[0] ;
 wire \osr.sample_count_r[1] ;
 wire \osr.sample_count_r[2] ;
 wire \osr.sample_count_r[3] ;
 wire \osr.sample_count_r[4] ;
 wire \osr.sample_count_r[5] ;
 wire \osr.sample_count_r[6] ;
 wire \osr.sample_count_r[7] ;
 wire \osr.sample_count_r[8] ;
 wire net3;
 wire net2;
 wire net1;

 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0627_ (.I(\cnb.sampled_avg_control_r[2] ),
    .ZN(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0628_ (.A1(\cnb.sampled_avg_control_r[1] ),
    .A2(\cnb.sampled_avg_control_r[0] ),
    .ZN(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _0629_ (.A1(_0167_),
    .A2(_0168_),
    .ZN(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0630_ (.I(net72),
    .ZN(net13));
 gf180mcu_fd_sc_mcu7t5v0__or3_4 _0631_ (.A1(\cnb.shift_register_r[4] ),
    .A2(\cnb.shift_register_r[5] ),
    .A3(\cnb.shift_register_r[6] ),
    .Z(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__or4_4 _0632_ (.A1(\cnb.shift_register_r[8] ),
    .A2(\cnb.shift_register_r[11] ),
    .A3(\cnb.shift_register_r[10] ),
    .A4(\cnb.shift_register_r[14] ),
    .Z(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _0633_ (.A1(\cnb.shift_register_r[7] ),
    .A2(\cnb.shift_register_r[9] ),
    .Z(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__or3_4 _0634_ (.A1(_0169_),
    .A2(_0170_),
    .A3(_0171_),
    .Z(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0635_ (.I(_0172_),
    .ZN(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__or4_4 _0636_ (.A1(\cnb.shift_register_r[3] ),
    .A2(\cnb.shift_register_r[2] ),
    .A3(\cnb.is_holding_result_w ),
    .A4(net139),
    .Z(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _0637_ (.A1(\cnb.shift_register_r[13] ),
    .A2(_0174_),
    .Z(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0638_ (.I(\cnb.shift_register_r[3] ),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _0639_ (.A1(\cnb.is_holding_result_w ),
    .A2(net139),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _0640_ (.A1(\cnb.is_holding_result_w ),
    .A2(net139),
    .Z(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__inv_8 _0641_ (.I(\cnb.shift_register_r[2] ),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0642_ (.I0(_0177_),
    .I1(_0178_),
    .S(_0179_),
    .Z(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output29 (.I(net29),
    .Z(a_nmatrix_col_out_n[0]));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _0644_ (.A1(\cnb.shift_register_r[3] ),
    .A2(_0179_),
    .A3(_0177_),
    .Z(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _0645_ (.A1(_0176_),
    .A2(_0180_),
    .B(_0182_),
    .C(\cnb.shift_register_r[13] ),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0646_ (.I(\cnb.shift_register_r[12] ),
    .ZN(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__or3_4 _0647_ (.A1(_0184_),
    .A2(\cnb.shift_register_r[13] ),
    .A3(_0174_),
    .Z(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _0648_ (.A1(\cnb.shift_register_r[12] ),
    .A2(_0175_),
    .A3(_0183_),
    .B(_0185_),
    .ZN(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _0649_ (.A1(\cnb.shift_register_r[12] ),
    .A2(\cnb.shift_register_r[13] ),
    .Z(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _0650_ (.A1(\cnb.shift_register_r[7] ),
    .A2(\cnb.shift_register_r[11] ),
    .A3(\cnb.shift_register_r[14] ),
    .Z(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__or4_4 _0651_ (.A1(_0169_),
    .A2(_0174_),
    .A3(_0187_),
    .A4(_0188_),
    .Z(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _0652_ (.A1(\cnb.shift_register_r[8] ),
    .A2(\cnb.shift_register_r[10] ),
    .ZN(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _0653_ (.A1(\cnb.shift_register_r[8] ),
    .A2(\cnb.shift_register_r[10] ),
    .Z(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0654_ (.I0(_0190_),
    .I1(_0191_),
    .S(\cnb.shift_register_r[9] ),
    .Z(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0655_ (.A1(_0189_),
    .A2(_0192_),
    .ZN(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0656_ (.A1(_0173_),
    .A2(_0186_),
    .B(_0193_),
    .ZN(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0657_ (.I(\cnb.shift_register_r[6] ),
    .ZN(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _0658_ (.A1(\cnb.shift_register_r[7] ),
    .A2(\cnb.shift_register_r[9] ),
    .ZN(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _0659_ (.A1(_0194_),
    .A2(_0195_),
    .Z(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _0660_ (.A1(\cnb.shift_register_r[6] ),
    .A2(_0171_),
    .Z(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _0661_ (.A1(_0170_),
    .A2(_0196_),
    .A3(_0197_),
    .Z(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _0662_ (.I(\cnb.shift_register_r[4] ),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _0663_ (.A1(_0199_),
    .A2(\cnb.shift_register_r[6] ),
    .A3(_0170_),
    .A4(_0171_),
    .Z(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0664_ (.A1(\cnb.shift_register_r[4] ),
    .A2(_0198_),
    .B(_0200_),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _0665_ (.A1(_0174_),
    .A2(_0187_),
    .Z(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0666_ (.A1(\cnb.shift_register_r[5] ),
    .A2(_0202_),
    .ZN(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _0667_ (.A1(\cnb.shift_register_r[7] ),
    .A2(\cnb.shift_register_r[14] ),
    .Z(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0668_ (.I(\cnb.shift_register_r[11] ),
    .ZN(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _0669_ (.A1(\cnb.shift_register_r[9] ),
    .A2(_0205_),
    .A3(_0191_),
    .Z(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__or4_4 _0670_ (.A1(_0169_),
    .A2(_0202_),
    .A3(_0204_),
    .A4(_0206_),
    .Z(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0671_ (.I(_0207_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0672_ (.A1(_0201_),
    .A2(_0203_),
    .B(_0208_),
    .ZN(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0673_ (.I(_0034_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0674_ (.I(net1),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__and3_4 _0675_ (.A1(_0176_),
    .A2(_0179_),
    .A3(_0199_),
    .Z(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _0676_ (.A1(_0020_),
    .A2(_0211_),
    .Z(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0677_ (.I(_0019_),
    .ZN(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0678_ (.A1(\cnb.average_counter_r[0] ),
    .A2(_0022_),
    .B(_0021_),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0679_ (.I(_0018_),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0680_ (.A1(_0213_),
    .A2(_0214_),
    .B(_0215_),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _0681_ (.A1(_0013_),
    .A2(_0016_),
    .Z(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _0682_ (.A1(_0013_),
    .A2(_0015_),
    .Z(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _0683_ (.A1(_0216_),
    .A2(_0217_),
    .B(_0218_),
    .C(_0012_),
    .ZN(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0684_ (.I0(\cnb.average_sum_r[2] ),
    .I1(\cnb.average_sum_r[3] ),
    .S(\cnb.sampled_avg_control_r[0] ),
    .Z(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0685_ (.A1(\cnb.sampled_avg_control_r[1] ),
    .A2(_0167_),
    .ZN(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0686_ (.A1(_0220_),
    .A2(_0221_),
    .ZN(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _0687_ (.A1(\cnb.sampled_avg_control_r[0] ),
    .A2(_0167_),
    .A3(\cnb.average_sum_r[4] ),
    .Z(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0688_ (.I(\cnb.sampled_avg_control_r[0] ),
    .ZN(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _0689_ (.A1(_0224_),
    .A2(\cnb.sampled_avg_control_r[2] ),
    .A3(\cnb.average_sum_r[1] ),
    .Z(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0690_ (.A1(_0223_),
    .A2(_0225_),
    .B(\cnb.sampled_avg_control_r[1] ),
    .ZN(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__or3_4 _0691_ (.A1(_0219_),
    .A2(_0222_),
    .A3(_0226_),
    .Z(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__or3_4 _0692_ (.A1(\cnb.shift_register_r[3] ),
    .A2(\cnb.shift_register_r[2] ),
    .A3(\cnb.shift_register_r[4] ),
    .Z(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _0693_ (.A1(_0210_),
    .A2(_0212_),
    .B1(_0227_),
    .B2(_0228_),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output28 (.I(net28),
    .Z(a_nmatrix_col_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0695_ (.I0(_0036_),
    .I1(_0209_),
    .S(_0229_),
    .Z(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0696_ (.I(_0004_),
    .ZN(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0697_ (.I(_0005_),
    .ZN(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _0698_ (.A1(_0184_),
    .A2(\cnb.shift_register_r[13] ),
    .A3(_0172_),
    .A4(_0174_),
    .Z(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _0699_ (.A1(\cnb.shift_register_r[9] ),
    .A2(\cnb.shift_register_r[8] ),
    .ZN(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _0700_ (.A1(\cnb.shift_register_r[10] ),
    .A2(_0189_),
    .A3(_0232_),
    .Z(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _0701_ (.A1(_0231_),
    .A2(_0233_),
    .Z(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0702_ (.I(\cnb.shift_register_r[10] ),
    .ZN(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__or4_4 _0703_ (.A1(\cnb.shift_register_r[9] ),
    .A2(\cnb.shift_register_r[8] ),
    .A3(_0235_),
    .A4(_0189_),
    .Z(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _0704_ (.A1(\cnb.shift_register_r[5] ),
    .A2(\cnb.shift_register_r[6] ),
    .Z(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0705_ (.A1(_0199_),
    .A2(_0237_),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _0706_ (.A1(_0170_),
    .A2(_0171_),
    .A3(_0202_),
    .A4(_0238_),
    .Z(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _0707_ (.A1(_0236_),
    .A2(_0239_),
    .Z(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _0708_ (.A1(\cnb.shift_register_r[12] ),
    .A2(\cnb.shift_register_r[13] ),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _0709_ (.A1(_0172_),
    .A2(_0174_),
    .A3(_0241_),
    .Z(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _0710_ (.A1(_0207_),
    .A2(_0242_),
    .Z(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _0711_ (.A1(_0169_),
    .A2(_0170_),
    .A3(_0202_),
    .A4(_0195_),
    .Z(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__and3_4 _0712_ (.A1(_0236_),
    .A2(_0243_),
    .A3(_0244_),
    .Z(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__and3_4 _0713_ (.A1(_0035_),
    .A2(_0240_),
    .A3(_0245_),
    .Z(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0714_ (.A1(_0234_),
    .A2(_0246_),
    .B(_0229_),
    .ZN(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _0715_ (.A1(\cnb.data_register_r[7] ),
    .A2(\cnb.data_register_r[8] ),
    .ZN(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__inv_8 _0716_ (.I(\cnb.data_register_r[9] ),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output27 (.I(net27),
    .Z(a_nmatrix_col_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__inv_8 _0718_ (.I(net8),
    .ZN(net52));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output26 (.I(net26),
    .Z(a_nmatrix_col_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _0720_ (.A1(_0248_),
    .A2(net52),
    .Z(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0721_ (.A1(_0247_),
    .A2(_0251_),
    .ZN(net42));
 gf180mcu_fd_sc_mcu7t5v0__inv_8 _0722_ (.I(\cnb.data_register_r[7] ),
    .ZN(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _0723_ (.A1(_0252_),
    .A2(\cnb.data_register_r[8] ),
    .Z(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0724_ (.A1(_0248_),
    .A2(_0253_),
    .ZN(net106));
 gf180mcu_fd_sc_mcu7t5v0__or3_4 _0725_ (.A1(net6),
    .A2(net5),
    .A3(net7),
    .Z(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0726_ (.I(_0082_),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _0727_ (.A1(\osr.sample_count_r[6] ),
    .A2(\osr.sample_count_r[8] ),
    .Z(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _0728_ (.A1(\osr.sample_count_r[3] ),
    .A2(\osr.sample_count_r[4] ),
    .A3(\osr.sample_count_r[5] ),
    .A4(\osr.sample_count_r[7] ),
    .Z(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__or4_4 _0729_ (.A1(\osr.sample_count_r[2] ),
    .A2(_0255_),
    .A3(_0256_),
    .A4(_0257_),
    .Z(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _0730_ (.A1(_0254_),
    .A2(_0258_),
    .Z(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output25 (.I(net25),
    .Z(a_nmatrix_col_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0732_ (.I(_0062_),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0733_ (.I(_0061_),
    .ZN(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0734_ (.I(_0067_),
    .ZN(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _0735_ (.A1(_0009_),
    .A2(_0261_),
    .B(_0262_),
    .C(_0263_),
    .ZN(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _0736_ (.A1(_0068_),
    .A2(_0067_),
    .B(_0072_),
    .C(_0066_),
    .ZN(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0737_ (.I(_0265_),
    .ZN(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0738_ (.A1(_0072_),
    .A2(_0065_),
    .B(_0071_),
    .ZN(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0739_ (.A1(_0069_),
    .A2(_0075_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0740_ (.A1(_0267_),
    .A2(_0268_),
    .ZN(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0741_ (.A1(_0264_),
    .A2(_0266_),
    .B(_0269_),
    .ZN(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0742_ (.I(_0075_),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0743_ (.A1(_0070_),
    .A2(_0069_),
    .B(_0076_),
    .ZN(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0744_ (.A1(_0271_),
    .A2(_0272_),
    .ZN(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _0745_ (.A1(_0074_),
    .A2(_0078_),
    .A3(_0273_),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0746_ (.A1(_0078_),
    .A2(_0073_),
    .B(_0077_),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0747_ (.A1(_0270_),
    .A2(_0274_),
    .B(_0275_),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _0748_ (.A1(\osr.result_r[10] ),
    .A2(_0276_),
    .Z(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _0749_ (.A1(_0259_),
    .A2(_0277_),
    .Z(\osr.next_result_w[10] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _0750_ (.A1(_0254_),
    .A2(_0258_),
    .ZN(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0751_ (.I(_0009_),
    .ZN(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _0752_ (.A1(_0279_),
    .A2(_0062_),
    .B(_0061_),
    .C(_0067_),
    .ZN(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _0753_ (.A1(_0280_),
    .A2(_0265_),
    .B(_0267_),
    .C(_0268_),
    .ZN(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__and3_4 _0754_ (.A1(_0074_),
    .A2(_0281_),
    .A3(_0273_),
    .Z(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0755_ (.A1(_0281_),
    .A2(_0273_),
    .B(_0074_),
    .ZN(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0756_ (.A1(\cnb.result_out[8] ),
    .A2(_0278_),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _0757_ (.A1(_0278_),
    .A2(_0282_),
    .A3(_0283_),
    .B(_0284_),
    .ZN(\osr.next_result_w[8] ));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0758_ (.A1(_0280_),
    .A2(_0265_),
    .B(_0267_),
    .ZN(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _0759_ (.A1(_0070_),
    .A2(_0285_),
    .Z(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0760_ (.I0(\cnb.result_out[6] ),
    .I1(_0286_),
    .S(_0259_),
    .Z(\osr.next_result_w[6] ));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0761_ (.A1(_0009_),
    .A2(_0261_),
    .B(_0262_),
    .ZN(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0762_ (.A1(_0068_),
    .A2(_0287_),
    .B(_0067_),
    .ZN(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _0763_ (.A1(_0066_),
    .A2(_0288_),
    .ZN(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0764_ (.I0(\cnb.result_out[4] ),
    .I1(_0289_),
    .S(_0259_),
    .Z(\osr.next_result_w[4] ));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _0765_ (.A1(_0079_),
    .A2(_0064_),
    .B(_0061_),
    .C(_0063_),
    .ZN(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0766_ (.A1(_0062_),
    .A2(_0061_),
    .B(_0068_),
    .ZN(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0767_ (.A1(_0065_),
    .A2(_0067_),
    .ZN(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0768_ (.A1(_0070_),
    .A2(_0071_),
    .B(_0069_),
    .ZN(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _0769_ (.A1(_0290_),
    .A2(_0291_),
    .B(_0292_),
    .C(_0293_),
    .ZN(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _0770_ (.A1(_0066_),
    .A2(_0065_),
    .B(_0072_),
    .C(_0070_),
    .ZN(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0771_ (.A1(_0074_),
    .A2(_0076_),
    .ZN(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0772_ (.A1(_0293_),
    .A2(_0295_),
    .B(_0296_),
    .ZN(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _0773_ (.A1(_0074_),
    .A2(_0075_),
    .Z(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _0774_ (.A1(_0073_),
    .A2(_0077_),
    .A3(_0298_),
    .Z(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0775_ (.A1(_0294_),
    .A2(_0297_),
    .B(_0299_),
    .ZN(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _0776_ (.A1(_0078_),
    .A2(_0077_),
    .Z(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0777_ (.A1(\osr.result_r[10] ),
    .A2(_0301_),
    .ZN(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0778_ (.A1(_0300_),
    .A2(_0302_),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _0779_ (.A1(\osr.result_r[11] ),
    .A2(_0303_),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0780_ (.A1(_0278_),
    .A2(_0304_),
    .ZN(\osr.next_result_w[11] ));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _0781_ (.A1(_0294_),
    .A2(_0297_),
    .B(_0298_),
    .C(_0073_),
    .ZN(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _0782_ (.A1(_0078_),
    .A2(_0305_),
    .ZN(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _0783_ (.A1(\cnb.result_out[9] ),
    .A2(_0278_),
    .Z(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0784_ (.A1(_0259_),
    .A2(_0306_),
    .B(_0307_),
    .ZN(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _0785_ (.I(_0308_),
    .ZN(\osr.next_result_w[9] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0786_ (.I(\cnb.result_out[7] ),
    .ZN(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0787_ (.A1(_0293_),
    .A2(_0295_),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _0788_ (.A1(_0294_),
    .A2(_0310_),
    .Z(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _0789_ (.A1(_0076_),
    .A2(_0311_),
    .ZN(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0790_ (.I0(_0309_),
    .I1(_0312_),
    .S(_0259_),
    .Z(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0791_ (.I(_0313_),
    .ZN(\osr.next_result_w[7] ));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0792_ (.A1(_0290_),
    .A2(_0291_),
    .B(_0263_),
    .ZN(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0793_ (.A1(_0066_),
    .A2(_0314_),
    .B(_0065_),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _0794_ (.A1(_0072_),
    .A2(_0315_),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0795_ (.I0(\cnb.result_out[5] ),
    .I1(_0316_),
    .S(_0259_),
    .Z(\osr.next_result_w[5] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output24 (.I(net24),
    .Z(a_nmatrix_col_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _0797_ (.A1(\osr.result_r[10] ),
    .A2(\osr.result_r[11] ),
    .A3(_0276_),
    .Z(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _0798_ (.A1(\osr.result_r[12] ),
    .A2(_0318_),
    .Z(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _0799_ (.A1(_0259_),
    .A2(_0319_),
    .Z(\osr.next_result_w[12] ));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _0800_ (.A1(\osr.result_r[10] ),
    .A2(\osr.result_r[11] ),
    .A3(\osr.result_r[12] ),
    .Z(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0801_ (.A1(_0301_),
    .A2(_0320_),
    .ZN(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _0802_ (.A1(_0300_),
    .A2(_0321_),
    .Z(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _0803_ (.A1(\osr.result_r[13] ),
    .A2(_0322_),
    .ZN(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _0804_ (.A1(_0259_),
    .A2(_0323_),
    .Z(\osr.next_result_w[13] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0805_ (.I(\osr.result_r[14] ),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _0806_ (.A1(\osr.result_r[13] ),
    .A2(_0320_),
    .Z(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _0807_ (.A1(_0276_),
    .A2(_0325_),
    .Z(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _0808_ (.A1(_0324_),
    .A2(_0326_),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _0809_ (.A1(_0259_),
    .A2(_0327_),
    .Z(\osr.next_result_w[14] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0810_ (.A1(_0301_),
    .A2(_0325_),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _0811_ (.A1(_0324_),
    .A2(_0300_),
    .A3(_0328_),
    .Z(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _0812_ (.A1(\osr.result_r[15] ),
    .A2(_0329_),
    .ZN(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _0813_ (.A1(_0259_),
    .A2(_0330_),
    .Z(\osr.next_result_w[15] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output23 (.I(net23),
    .Z(a_nmatrix_col_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _0815_ (.A1(\cnb.data_register_r[9] ),
    .A2(net52),
    .Z(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _0816_ (.A1(\cnb.data_register_r[7] ),
    .A2(\cnb.data_register_r[8] ),
    .Z(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0817_ (.A1(_0332_),
    .A2(_0333_),
    .ZN(net101));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _0818_ (.I(\cnb.data_register_r[8] ),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _0819_ (.A1(\cnb.data_register_r[7] ),
    .A2(_0334_),
    .Z(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0820_ (.A1(\cnb.data_register_r[9] ),
    .A2(_0335_),
    .ZN(net47));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0821_ (.I(\cnb.result_out[1] ),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0822_ (.I(\osr.result_r[1] ),
    .ZN(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0823_ (.I(_0079_),
    .ZN(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0824_ (.A1(\cnb.sampled_avg_control_r[2] ),
    .A2(_0168_),
    .ZN(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0825_ (.I(_0221_),
    .ZN(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _0826_ (.A1(\cnb.sampled_avg_control_r[2] ),
    .A2(_0168_),
    .B1(_0336_),
    .B2(\cnb.sampled_avg_control_r[0] ),
    .ZN(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _0827_ (.A1(_0221_),
    .A2(_0011_),
    .Z(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _0828_ (.A1(_0033_),
    .A2(_0034_),
    .A3(_0240_),
    .Z(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0829_ (.A1(_0229_),
    .A2(_0337_),
    .ZN(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0830_ (.I(\cnb.shift_register_r[13] ),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _0831_ (.A1(\cnb.shift_register_r[12] ),
    .A2(_0339_),
    .A3(_0172_),
    .A4(_0174_),
    .Z(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0832_ (.I0(_0229_),
    .I1(_0338_),
    .S(_0340_),
    .Z(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _0833_ (.I(net73),
    .ZN(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0834_ (.I(_0033_),
    .ZN(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0835_ (.A1(_0035_),
    .A2(_0229_),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _0836_ (.A1(_0240_),
    .A2(_0341_),
    .ZN(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _0837_ (.A1(_0245_),
    .A2(_0338_),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0838_ (.A1(_0229_),
    .A2(_0246_),
    .ZN(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _0839_ (.A1(_0234_),
    .A2(_0342_),
    .ZN(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _0840_ (.A1(_0231_),
    .A2(_0236_),
    .Z(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _0841_ (.A1(_0338_),
    .A2(_0343_),
    .ZN(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0842_ (.I0(_0229_),
    .I1(_0058_),
    .S(_0243_),
    .Z(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0843_ (.I(\osr.sample_count_r[1] ),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _0844_ (.A1(_0179_),
    .A2(_0032_),
    .Z(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _0845_ (.A1(_0216_),
    .A2(_0217_),
    .Z(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__or3_4 _0846_ (.A1(_0012_),
    .A2(_0345_),
    .A3(_0218_),
    .Z(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _0847_ (.A1(_0211_),
    .A2(_0346_),
    .Z(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output22 (.I(net22),
    .Z(a_nmatrix_col_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0849_ (.I0(net72),
    .I1(_0344_),
    .S(_0347_),
    .Z(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _0850_ (.A1(_0177_),
    .A2(_0349_),
    .Z(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0851_ (.A1(\cnb.shift_register_r[2] ),
    .A2(_0003_),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0852_ (.I0(net73),
    .I1(_0350_),
    .S(_0347_),
    .Z(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _0853_ (.A1(_0177_),
    .A2(_0351_),
    .Z(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _0854_ (.A1(_0002_),
    .A2(_0041_),
    .ZN(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _0855_ (.A1(_0179_),
    .A2(_0352_),
    .Z(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0856_ (.I0(net74),
    .I1(_0353_),
    .S(_0347_),
    .Z(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _0857_ (.A1(_0177_),
    .A2(_0354_),
    .Z(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output21 (.I(net21),
    .Z(a_nmatrix_col_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0859_ (.I(_0041_),
    .ZN(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0860_ (.A1(_0005_),
    .A2(_0038_),
    .B(_0037_),
    .ZN(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0861_ (.A1(_0356_),
    .A2(_0357_),
    .ZN(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _0862_ (.A1(_0044_),
    .A2(_0040_),
    .A3(_0358_),
    .Z(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _0863_ (.A1(_0005_),
    .A2(_0038_),
    .B(_0037_),
    .C(_0040_),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0864_ (.A1(_0041_),
    .A2(_0040_),
    .B(_0044_),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _0865_ (.A1(_0360_),
    .A2(_0361_),
    .Z(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _0866_ (.A1(_0179_),
    .A2(_0359_),
    .A3(_0362_),
    .Z(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0867_ (.I0(\cnb.data_register_r[3] ),
    .I1(_0363_),
    .S(_0347_),
    .Z(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _0868_ (.A1(_0177_),
    .A2(_0364_),
    .Z(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output20 (.I(net20),
    .Z(a_nmatrix_col_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0870_ (.I(_0040_),
    .ZN(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0871_ (.A1(_0002_),
    .A2(_0356_),
    .B(_0366_),
    .ZN(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0872_ (.A1(_0044_),
    .A2(_0367_),
    .B(_0043_),
    .ZN(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _0873_ (.A1(_0047_),
    .A2(_0368_),
    .ZN(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _0874_ (.A1(_0179_),
    .A2(_0369_),
    .Z(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0875_ (.I0(\cnb.data_register_r[4] ),
    .I1(_0370_),
    .S(_0347_),
    .Z(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _0876_ (.A1(_0177_),
    .A2(_0371_),
    .Z(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output19 (.I(net19),
    .Z(a_nmatrix_col_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _0878_ (.A1(_0211_),
    .A2(_0346_),
    .ZN(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output18 (.I(net18),
    .Z(a_nmatrix_col_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output17 (.I(net17),
    .Z(a_nmatrix_col_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0881_ (.A1(\cnb.data_register_r[5] ),
    .A2(_0373_),
    .ZN(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0882_ (.I(_0046_),
    .ZN(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0883_ (.A1(_0360_),
    .A2(_0361_),
    .ZN(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0884_ (.A1(_0043_),
    .A2(_0378_),
    .B(_0047_),
    .ZN(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _0885_ (.A1(_0050_),
    .A2(_0377_),
    .A3(_0379_),
    .Z(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0886_ (.A1(_0377_),
    .A2(_0379_),
    .B(_0050_),
    .ZN(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output16 (.I(net16),
    .Z(a_nmatrix_col_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _0888_ (.A1(_0380_),
    .A2(_0381_),
    .B(_0179_),
    .C(_0347_),
    .ZN(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _0889_ (.A1(\cnb.is_holding_result_w ),
    .A2(net139),
    .Z(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0890_ (.A1(_0376_),
    .A2(_0383_),
    .B(_0384_),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output15 (.I(net15),
    .Z(a_nmatrix_bincap_out_n[2]));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0892_ (.A1(\cnb.data_register_r[6] ),
    .A2(_0373_),
    .ZN(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0893_ (.I(_0047_),
    .ZN(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0894_ (.A1(_0387_),
    .A2(_0368_),
    .B(_0377_),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0895_ (.A1(_0050_),
    .A2(_0388_),
    .B(_0049_),
    .ZN(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _0896_ (.A1(_0053_),
    .A2(_0389_),
    .Z(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _0897_ (.A1(\cnb.shift_register_r[2] ),
    .A2(_0373_),
    .A3(_0390_),
    .Z(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0898_ (.A1(_0386_),
    .A2(_0391_),
    .B(_0384_),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _0899_ (.A1(_0053_),
    .A2(_0049_),
    .Z(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _0900_ (.A1(_0043_),
    .A2(_0046_),
    .A3(_0052_),
    .A4(_0392_),
    .ZN(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _0901_ (.A1(_0050_),
    .A2(_0057_),
    .Z(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _0902_ (.A1(_0047_),
    .A2(_0046_),
    .Z(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _0903_ (.A1(_0394_),
    .A2(_0395_),
    .B(_0052_),
    .C(_0392_),
    .ZN(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0904_ (.A1(_0362_),
    .A2(_0393_),
    .B(_0396_),
    .ZN(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _0905_ (.A1(_0056_),
    .A2(_0397_),
    .Z(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _0906_ (.A1(_0179_),
    .A2(_0398_),
    .Z(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0907_ (.I0(\cnb.data_register_r[7] ),
    .I1(_0399_),
    .S(_0347_),
    .Z(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _0908_ (.A1(_0177_),
    .A2(_0400_),
    .Z(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _0909_ (.A1(_0179_),
    .A2(_0060_),
    .A3(_0177_),
    .A4(_0347_),
    .ZN(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _0910_ (.A1(\cnb.shift_register_r[2] ),
    .A2(_0060_),
    .A3(_0384_),
    .A4(_0373_),
    .Z(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0911_ (.A1(_0053_),
    .A2(_0056_),
    .ZN(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0912_ (.A1(_0056_),
    .A2(_0052_),
    .B(_0055_),
    .ZN(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0913_ (.A1(_0389_),
    .A2(_0403_),
    .B(_0404_),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0914_ (.I0(_0401_),
    .I1(_0402_),
    .S(_0405_),
    .Z(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _0915_ (.A1(_0334_),
    .A2(_0384_),
    .A3(_0347_),
    .B(_0406_),
    .ZN(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _0916_ (.A1(_0056_),
    .A2(_0060_),
    .A3(_0397_),
    .Z(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _0917_ (.A1(_0060_),
    .A2(_0055_),
    .B(_0059_),
    .C(_0407_),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0918_ (.A1(_0179_),
    .A2(\cnb.data_register_r[9] ),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _0919_ (.A1(_0384_),
    .A2(_0373_),
    .A3(_0408_),
    .A4(_0409_),
    .Z(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _0920_ (.A1(\cnb.shift_register_r[2] ),
    .A2(\cnb.data_register_r[9] ),
    .A3(_0384_),
    .A4(_0408_),
    .Z(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0921_ (.A1(_0172_),
    .A2(_0185_),
    .ZN(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _0922_ (.A1(\cnb.shift_register_r[12] ),
    .A2(_0172_),
    .A3(_0175_),
    .A4(_0183_),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _0923_ (.A1(_0193_),
    .A2(_0412_),
    .A3(_0413_),
    .ZN(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _0924_ (.A1(\cnb.shift_register_r[4] ),
    .A2(\cnb.shift_register_r[5] ),
    .A3(_0202_),
    .A4(_0198_),
    .Z(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _0925_ (.A1(\cnb.shift_register_r[9] ),
    .A2(_0205_),
    .A3(_0169_),
    .A4(_0204_),
    .Z(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _0926_ (.A1(_0191_),
    .A2(_0174_),
    .A3(_0187_),
    .A4(_0416_),
    .Z(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _0927_ (.A1(\cnb.shift_register_r[5] ),
    .A2(_0202_),
    .A3(_0200_),
    .Z(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _0928_ (.A1(_0415_),
    .A2(_0417_),
    .A3(_0418_),
    .A4(_0240_),
    .Z(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0929_ (.A1(_0414_),
    .A2(_0419_),
    .B(_0229_),
    .ZN(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0930_ (.I0(_0410_),
    .I1(_0411_),
    .S(_0420_),
    .Z(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _0931_ (.A1(_0179_),
    .A2(_0248_),
    .A3(_0177_),
    .A4(_0408_),
    .ZN(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0932_ (.A1(_0384_),
    .A2(_0409_),
    .ZN(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _0933_ (.A1(_0347_),
    .A2(_0408_),
    .A3(_0423_),
    .ZN(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0934_ (.I0(_0422_),
    .I1(_0424_),
    .S(_0420_),
    .Z(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _0935_ (.A1(\cnb.data_register_r[9] ),
    .A2(_0384_),
    .A3(_0347_),
    .Z(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _0936_ (.A1(_0421_),
    .A2(_0425_),
    .A3(_0426_),
    .Z(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _0937_ (.A1(net72),
    .A2(_0229_),
    .ZN(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _0938_ (.A1(\cnb.shift_register_r[2] ),
    .A2(_0346_),
    .Z(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output14 (.I(net14),
    .Z(a_nmatrix_bincap_out_n[1]));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0940_ (.I0(\cnb.result_out[0] ),
    .I1(_0427_),
    .S(_0428_),
    .Z(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0941_ (.I(_0030_),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0942_ (.I0(_0430_),
    .I1(net73),
    .S(_0229_),
    .Z(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0943_ (.I0(\cnb.result_out[1] ),
    .I1(_0431_),
    .S(_0428_),
    .Z(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0944_ (.I(net74),
    .ZN(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0945_ (.I(_0029_),
    .ZN(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0946_ (.A1(_0432_),
    .A2(_0229_),
    .ZN(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _0947_ (.A1(net15),
    .A2(_0433_),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0948_ (.I0(\cnb.result_out[2] ),
    .I1(_0434_),
    .S(_0428_),
    .Z(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0949_ (.I(\cnb.data_register_r[3] ),
    .ZN(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__or3_4 _0950_ (.A1(net73),
    .A2(net74),
    .A3(net72),
    .Z(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0951_ (.A1(_0229_),
    .A2(_0436_),
    .ZN(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _0952_ (.A1(_0435_),
    .A2(_0437_),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0953_ (.I0(\cnb.result_out[3] ),
    .I1(_0438_),
    .S(_0428_),
    .Z(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _0954_ (.A1(_0432_),
    .A2(net74),
    .A3(\cnb.data_register_r[3] ),
    .A4(_0229_),
    .Z(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _0955_ (.A1(\cnb.data_register_r[4] ),
    .A2(_0439_),
    .ZN(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0956_ (.I0(\cnb.result_out[4] ),
    .I1(_0440_),
    .S(_0428_),
    .Z(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _0957_ (.A1(\cnb.data_register_r[3] ),
    .A2(\cnb.data_register_r[4] ),
    .A3(_0229_),
    .A4(_0436_),
    .Z(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _0958_ (.A1(\cnb.data_register_r[5] ),
    .A2(_0441_),
    .ZN(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0959_ (.I0(\cnb.result_out[5] ),
    .I1(_0442_),
    .S(_0428_),
    .Z(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__or3_4 _0960_ (.A1(\cnb.data_register_r[3] ),
    .A2(\cnb.data_register_r[4] ),
    .A3(\cnb.data_register_r[5] ),
    .Z(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _0961_ (.A1(_0432_),
    .A2(net74),
    .A3(_0229_),
    .A4(_0443_),
    .Z(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _0962_ (.A1(\cnb.data_register_r[6] ),
    .A2(_0444_),
    .ZN(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0963_ (.I0(\cnb.result_out[6] ),
    .I1(_0445_),
    .S(_0428_),
    .Z(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _0964_ (.A1(\cnb.data_register_r[6] ),
    .A2(_0443_),
    .Z(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _0965_ (.A1(_0229_),
    .A2(_0436_),
    .A3(_0446_),
    .Z(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _0966_ (.A1(\cnb.data_register_r[7] ),
    .A2(_0447_),
    .ZN(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0967_ (.I0(\cnb.result_out[7] ),
    .I1(_0448_),
    .S(_0428_),
    .Z(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0968_ (.A1(\cnb.data_register_r[6] ),
    .A2(_0443_),
    .ZN(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0969_ (.A1(_0252_),
    .A2(_0449_),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _0970_ (.A1(_0432_),
    .A2(net74),
    .A3(_0229_),
    .A4(_0450_),
    .Z(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _0971_ (.A1(\cnb.data_register_r[8] ),
    .A2(_0451_),
    .ZN(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0972_ (.I0(\cnb.result_out[8] ),
    .I1(_0452_),
    .S(_0428_),
    .Z(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0973_ (.A1(_0252_),
    .A2(_0334_),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _0974_ (.A1(_0229_),
    .A2(_0453_),
    .A3(_0436_),
    .A4(_0446_),
    .Z(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _0975_ (.A1(\cnb.data_register_r[9] ),
    .A2(_0454_),
    .ZN(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0976_ (.I0(\cnb.result_out[9] ),
    .I1(_0455_),
    .S(_0428_),
    .Z(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0977_ (.I0(\cnb.sampled_avg_control_r[0] ),
    .I1(net2),
    .S(net139),
    .Z(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0978_ (.I0(\cnb.sampled_avg_control_r[1] ),
    .I1(net3),
    .S(net139),
    .Z(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0979_ (.I0(\cnb.sampled_avg_control_r[2] ),
    .I1(net4),
    .S(net139),
    .Z(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0980_ (.I(_0258_),
    .ZN(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _0981_ (.A1(\osr.osr_mode_r[0] ),
    .A2(_0259_),
    .Z(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0982_ (.A1(net5),
    .A2(_0456_),
    .B(_0457_),
    .ZN(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0983_ (.I(_0458_),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output13 (.I(net13),
    .Z(a_nmatrix_bincap_out_n[0]));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0985_ (.I0(net6),
    .I1(\osr.osr_mode_r[1] ),
    .S(_0259_),
    .Z(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _0986_ (.A1(net7),
    .A2(_0456_),
    .B1(_0259_),
    .B2(\osr.osr_mode_r[2] ),
    .ZN(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0987_ (.I(_0460_),
    .ZN(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _0988_ (.A1(net131),
    .A2(_0254_),
    .Z(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__inv_8 _0989_ (.I(\osr.osr_mode_r[2] ),
    .ZN(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _0990_ (.I(\osr.osr_mode_r[0] ),
    .ZN(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _0991_ (.A1(_0009_),
    .A2(_0062_),
    .ZN(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _0992_ (.I0(\cnb.result_out[2] ),
    .I1(\cnb.result_out[6] ),
    .I2(_0464_),
    .I3(_0286_),
    .S0(\osr.osr_mode_r[1] ),
    .S1(_0259_),
    .Z(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0993_ (.A1(_0463_),
    .A2(\osr.osr_mode_r[1] ),
    .ZN(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _0994_ (.A1(_0463_),
    .A2(_0465_),
    .B1(_0466_),
    .B2(\osr.next_result_w[4] ),
    .ZN(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _0995_ (.A1(\osr.osr_mode_r[0] ),
    .A2(\osr.osr_mode_r[1] ),
    .ZN(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _0996_ (.A1(\osr.osr_mode_r[2] ),
    .A2(_0468_),
    .ZN(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0997_ (.A1(\osr.next_result_w[8] ),
    .A2(_0469_),
    .ZN(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0998_ (.A1(_0462_),
    .A2(_0467_),
    .B(_0470_),
    .ZN(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0999_ (.I(\osr.sample_count_r[6] ),
    .ZN(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _1000_ (.A1(\osr.osr_mode_r[1] ),
    .A2(\osr.osr_mode_r[2] ),
    .B1(\osr.sample_count_r[2] ),
    .B2(_0472_),
    .ZN(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _1001_ (.A1(\osr.osr_mode_r[1] ),
    .A2(_0462_),
    .ZN(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1002_ (.I(\osr.sample_count_r[2] ),
    .ZN(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1003_ (.A1(\osr.osr_mode_r[0] ),
    .A2(_0473_),
    .B1(_0474_),
    .B2(_0475_),
    .ZN(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _1004_ (.A1(\osr.osr_mode_r[0] ),
    .A2(\osr.sample_count_r[2] ),
    .A3(_0474_),
    .Z(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1005_ (.I0(_0476_),
    .I1(_0477_),
    .S(\osr.sample_count_r[4] ),
    .Z(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1006_ (.A1(\osr.sample_count_r[8] ),
    .A2(_0468_),
    .ZN(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _1007_ (.A1(\osr.sample_count_r[8] ),
    .A2(_0468_),
    .Z(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1008_ (.I0(_0479_),
    .I1(_0480_),
    .S(\osr.sample_count_r[0] ),
    .Z(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1009_ (.A1(\osr.sample_count_r[0] ),
    .A2(_0468_),
    .Z(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _1010_ (.A1(\osr.sample_count_r[8] ),
    .A2(_0482_),
    .Z(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1011_ (.I0(_0481_),
    .I1(_0483_),
    .S(_0462_),
    .Z(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _1012_ (.A1(_0463_),
    .A2(\osr.osr_mode_r[2] ),
    .A3(\osr.sample_count_r[2] ),
    .Z(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__and3_4 _1013_ (.A1(\osr.osr_mode_r[0] ),
    .A2(\osr.osr_mode_r[1] ),
    .A3(_0462_),
    .Z(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1014_ (.A1(_0472_),
    .A2(_0485_),
    .B(_0486_),
    .ZN(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _1015_ (.A1(\osr.sample_count_r[1] ),
    .A2(\osr.sample_count_r[3] ),
    .A3(\osr.sample_count_r[5] ),
    .A4(\osr.sample_count_r[7] ),
    .Z(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _1016_ (.A1(_0487_),
    .A2(_0488_),
    .Z(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1017_ (.A1(_0278_),
    .A2(_0478_),
    .A3(_0484_),
    .A4(_0489_),
    .ZN(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1018_ (.I0(_0461_),
    .I1(_0471_),
    .S(_0490_),
    .Z(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _1019_ (.A1(\osr.osr_mode_r[1] ),
    .A2(\osr.next_result_w[9] ),
    .B1(\osr.next_result_w[5] ),
    .B2(_0474_),
    .ZN(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1020_ (.A1(_0463_),
    .A2(_0491_),
    .Z(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1021_ (.A1(_0079_),
    .A2(_0064_),
    .B(_0063_),
    .ZN(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1022_ (.A1(_0261_),
    .A2(_0493_),
    .B(_0262_),
    .ZN(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1023_ (.A1(_0068_),
    .A2(_0494_),
    .Z(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1024_ (.I0(\cnb.result_out[3] ),
    .I1(_0495_),
    .S(_0259_),
    .Z(\osr.next_result_w[3] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1025_ (.A1(\osr.osr_mode_r[0] ),
    .A2(_0462_),
    .ZN(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _1026_ (.A1(\osr.osr_mode_r[1] ),
    .A2(_0496_),
    .Z(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _1027_ (.A1(\osr.next_result_w[3] ),
    .A2(_0497_),
    .Z(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1028_ (.A1(_0313_),
    .A2(_0486_),
    .ZN(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1029_ (.A1(\osr.osr_mode_r[2] ),
    .A2(_0308_),
    .ZN(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _1030_ (.A1(_0490_),
    .A2(_0498_),
    .A3(_0499_),
    .A4(_0500_),
    .ZN(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__or4_4 _1031_ (.A1(_0278_),
    .A2(_0478_),
    .A3(_0484_),
    .A4(_0489_),
    .Z(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _1032_ (.A1(_0254_),
    .A2(_0502_),
    .Z(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output12 (.I(net12),
    .Z(a_enable_loop_out));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1034_ (.A1(net132),
    .A2(_0503_),
    .ZN(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1035_ (.A1(_0492_),
    .A2(_0501_),
    .B(_0505_),
    .ZN(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1036_ (.A1(\osr.osr_mode_r[1] ),
    .A2(_0462_),
    .Z(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1037_ (.I0(\osr.next_result_w[8] ),
    .I1(\osr.next_result_w[6] ),
    .S(_0463_),
    .Z(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1038_ (.A1(_0506_),
    .A2(_0507_),
    .ZN(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1039_ (.A1(\osr.osr_mode_r[1] ),
    .A2(_0496_),
    .ZN(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1040_ (.A1(\osr.next_result_w[10] ),
    .A2(_0474_),
    .B(_0502_),
    .C(_0509_),
    .ZN(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1041_ (.A1(net133),
    .A2(_0254_),
    .ZN(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1042_ (.A1(\osr.next_result_w[4] ),
    .A2(_0497_),
    .ZN(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1043_ (.I0(_0511_),
    .I1(_0512_),
    .S(_0490_),
    .Z(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1044_ (.A1(_0508_),
    .A2(_0510_),
    .B(_0513_),
    .ZN(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1045_ (.A1(_0462_),
    .A2(_0313_),
    .ZN(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1046_ (.A1(\osr.osr_mode_r[1] ),
    .A2(_0278_),
    .A3(_0304_),
    .ZN(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1047_ (.A1(\osr.osr_mode_r[1] ),
    .A2(_0514_),
    .B(_0515_),
    .C(\osr.osr_mode_r[0] ),
    .ZN(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1048_ (.A1(_0308_),
    .A2(_0486_),
    .B(_0502_),
    .ZN(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _1049_ (.A1(_0462_),
    .A2(\osr.next_result_w[11] ),
    .B1(\osr.next_result_w[5] ),
    .B2(_0497_),
    .C(_0517_),
    .ZN(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1050_ (.A1(net134),
    .A2(_0503_),
    .ZN(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1051_ (.A1(_0516_),
    .A2(_0518_),
    .B(_0519_),
    .ZN(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1052_ (.A1(\osr.result_r[12] ),
    .A2(_0259_),
    .Z(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1053_ (.A1(\osr.result_r[10] ),
    .A2(\osr.result_r[11] ),
    .ZN(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1054_ (.A1(\osr.result_r[12] ),
    .A2(_0278_),
    .A3(_0521_),
    .ZN(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1055_ (.I0(_0520_),
    .I1(_0522_),
    .S(_0276_),
    .Z(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _1056_ (.A1(\osr.result_r[12] ),
    .A2(_0259_),
    .A3(_0521_),
    .Z(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _1057_ (.A1(\osr.osr_mode_r[1] ),
    .A2(_0523_),
    .A3(_0524_),
    .Z(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _1058_ (.A1(\osr.next_result_w[8] ),
    .A2(_0474_),
    .Z(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1059_ (.A1(_0525_),
    .A2(_0526_),
    .B(\osr.osr_mode_r[0] ),
    .ZN(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1060_ (.I0(\osr.next_result_w[6] ),
    .I1(_0277_),
    .S(\osr.osr_mode_r[1] ),
    .Z(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _1061_ (.A1(_0462_),
    .A2(_0319_),
    .B1(_0496_),
    .B2(_0528_),
    .C(_0490_),
    .ZN(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1062_ (.I(\cnb.result_out[0] ),
    .ZN(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1063_ (.A1(net135),
    .A2(_0502_),
    .ZN(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1064_ (.I0(_0530_),
    .I1(_0531_),
    .S(_0254_),
    .Z(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1065_ (.A1(_0527_),
    .A2(_0529_),
    .B(_0532_),
    .ZN(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1066_ (.I(_0469_),
    .ZN(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1067_ (.A1(\osr.next_result_w[11] ),
    .A2(_0486_),
    .B1(_0533_),
    .B2(\osr.next_result_w[13] ),
    .ZN(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1068_ (.A1(_0463_),
    .A2(_0506_),
    .Z(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _1069_ (.A1(\osr.next_result_w[7] ),
    .A2(_0509_),
    .B1(_0535_),
    .B2(\osr.next_result_w[9] ),
    .C(_0502_),
    .ZN(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1070_ (.A1(net136),
    .A2(_0490_),
    .ZN(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1071_ (.I0(_0006_),
    .I1(_0537_),
    .S(_0254_),
    .Z(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1072_ (.A1(_0534_),
    .A2(_0536_),
    .B(_0538_),
    .ZN(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1073_ (.A1(\osr.next_result_w[8] ),
    .A2(_0497_),
    .B(_0490_),
    .ZN(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1074_ (.A1(_0259_),
    .A2(_0327_),
    .B(_0469_),
    .ZN(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _1075_ (.A1(_0463_),
    .A2(\osr.next_result_w[10] ),
    .B1(_0319_),
    .B2(_0457_),
    .C(_0474_),
    .ZN(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1076_ (.I0(\cnb.result_out[2] ),
    .I1(net137),
    .S(_0254_),
    .Z(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1077_ (.A1(_0502_),
    .A2(_0542_),
    .ZN(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _1078_ (.A1(_0539_),
    .A2(_0540_),
    .A3(_0541_),
    .B(_0543_),
    .ZN(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1079_ (.I(\osr.result_r[13] ),
    .ZN(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1080_ (.A1(_0544_),
    .A2(_0322_),
    .Z(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1081_ (.I0(_0304_),
    .I1(_0545_),
    .S(\osr.osr_mode_r[0] ),
    .Z(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1082_ (.A1(_0300_),
    .A2(_0328_),
    .ZN(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _1083_ (.A1(_0278_),
    .A2(_0547_),
    .A3(_0474_),
    .A4(_0502_),
    .Z(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1084_ (.I(\cnb.result_out[3] ),
    .ZN(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1085_ (.A1(_0549_),
    .A2(_0254_),
    .ZN(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _1086_ (.A1(\osr.next_result_w[9] ),
    .A2(_0490_),
    .A3(_0509_),
    .Z(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1087_ (.A1(net138),
    .A2(_0503_),
    .B(_0550_),
    .C(_0551_),
    .ZN(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1088_ (.A1(\osr.next_result_w[15] ),
    .A2(_0490_),
    .A3(_0533_),
    .ZN(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1089_ (.A1(_0546_),
    .A2(_0548_),
    .B(_0552_),
    .C(_0553_),
    .ZN(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1090_ (.I0(\cnb.is_holding_result_w ),
    .I1(net139),
    .S(_0373_),
    .Z(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1091_ (.I0(\cnb.shift_register_r[11] ),
    .I1(\cnb.shift_register_r[10] ),
    .S(_0373_),
    .Z(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1092_ (.I0(\cnb.shift_register_r[11] ),
    .I1(\cnb.shift_register_r[12] ),
    .S(_0347_),
    .Z(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1093_ (.I0(\cnb.shift_register_r[12] ),
    .I1(\cnb.shift_register_r[13] ),
    .S(_0347_),
    .Z(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1094_ (.I0(\cnb.shift_register_r[13] ),
    .I1(\cnb.shift_register_r[14] ),
    .S(_0347_),
    .Z(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1095_ (.I0(net139),
    .I1(\cnb.shift_register_r[14] ),
    .S(_0373_),
    .Z(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1096_ (.A1(\cnb.is_holding_result_w ),
    .A2(_0373_),
    .Z(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _1097_ (.A1(_0428_),
    .A2(_0554_),
    .Z(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1098_ (.I0(\cnb.shift_register_r[3] ),
    .I1(\cnb.shift_register_r[2] ),
    .S(_0219_),
    .Z(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1099_ (.I0(\cnb.shift_register_r[4] ),
    .I1(\cnb.shift_register_r[3] ),
    .S(_0219_),
    .Z(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1100_ (.A1(\cnb.shift_register_r[5] ),
    .A2(_0347_),
    .ZN(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1101_ (.A1(_0199_),
    .A2(_0346_),
    .B(_0555_),
    .ZN(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1102_ (.I0(\cnb.shift_register_r[5] ),
    .I1(\cnb.shift_register_r[6] ),
    .S(_0347_),
    .Z(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1103_ (.I0(\cnb.shift_register_r[7] ),
    .I1(\cnb.shift_register_r[6] ),
    .S(_0373_),
    .Z(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1104_ (.I0(\cnb.shift_register_r[7] ),
    .I1(\cnb.shift_register_r[8] ),
    .S(_0347_),
    .Z(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1105_ (.I0(\cnb.shift_register_r[9] ),
    .I1(\cnb.shift_register_r[8] ),
    .S(_0373_),
    .Z(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1106_ (.I0(\cnb.shift_register_r[9] ),
    .I1(\cnb.shift_register_r[10] ),
    .S(_0347_),
    .Z(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1107_ (.A1(\cnb.conv_finished_r ),
    .A2(\osr.data_valid_r ),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1108_ (.I(net139),
    .ZN(net12));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _1109_ (.A1(_0248_),
    .A2(_0247_),
    .Z(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1110_ (.A1(net9),
    .A2(_0556_),
    .B(net8),
    .ZN(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__inv_8 _1111_ (.I(net9),
    .ZN(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _1112_ (.A1(_0252_),
    .A2(_0558_),
    .Z(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1113_ (.A1(_0446_),
    .A2(_0557_),
    .B(_0559_),
    .ZN(net29));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1114_ (.I(net29),
    .ZN(net16));
 gf180mcu_fd_sc_mcu7t5v0__inv_8 _1115_ (.I(\cnb.data_register_r[5] ),
    .ZN(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _1116_ (.A1(_0558_),
    .A2(net52),
    .Z(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output11 (.I(net11),
    .Z(a_conv_finished_osr_out));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _1118_ (.A1(_0248_),
    .A2(_0247_),
    .ZN(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _1119_ (.A1(net52),
    .A2(_0563_),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1120_ (.I(net53),
    .ZN(net62));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1121_ (.A1(net9),
    .A2(net62),
    .B(_0435_),
    .ZN(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1122_ (.A1(_0561_),
    .A2(_0564_),
    .B(\cnb.data_register_r[4] ),
    .ZN(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1123_ (.A1(_0560_),
    .A2(_0565_),
    .ZN(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _1124_ (.A1(\cnb.data_register_r[7] ),
    .A2(_0558_),
    .ZN(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _1125_ (.A1(\cnb.data_register_r[6] ),
    .A2(_0566_),
    .A3(_0567_),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _1126_ (.A1(\cnb.data_register_r[3] ),
    .A2(\cnb.data_register_r[4] ),
    .Z(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1127_ (.A1(_0568_),
    .A2(_0557_),
    .ZN(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _1128_ (.A1(\cnb.data_register_r[3] ),
    .A2(_0557_),
    .Z(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _1129_ (.A1(\cnb.data_register_r[4] ),
    .A2(_0570_),
    .Z(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1130_ (.A1(net9),
    .A2(_0571_),
    .ZN(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1131_ (.A1(net9),
    .A2(_0569_),
    .B(_0572_),
    .C(_0560_),
    .ZN(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _1132_ (.A1(\cnb.data_register_r[6] ),
    .A2(_0567_),
    .A3(_0573_),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__or3_4 _1133_ (.A1(\cnb.data_register_r[3] ),
    .A2(\cnb.data_register_r[4] ),
    .A3(_0557_),
    .Z(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1134_ (.A1(\cnb.data_register_r[6] ),
    .A2(_0252_),
    .A3(_0574_),
    .ZN(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1135_ (.A1(_0558_),
    .A2(_0569_),
    .B(_0575_),
    .ZN(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1136_ (.A1(\cnb.data_register_r[6] ),
    .A2(net9),
    .B1(_0576_),
    .B2(\cnb.data_register_r[5] ),
    .ZN(net32));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1137_ (.I(net32),
    .ZN(net19));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _1138_ (.I(\cnb.data_register_r[6] ),
    .ZN(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _1139_ (.A1(_0560_),
    .A2(_0577_),
    .Z(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1140_ (.A1(\cnb.data_register_r[4] ),
    .A2(_0570_),
    .ZN(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1141_ (.A1(_0578_),
    .A2(_0579_),
    .ZN(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1142_ (.A1(_0559_),
    .A2(_0580_),
    .ZN(net33));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1143_ (.I(net33),
    .ZN(net20));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1144_ (.A1(\cnb.data_register_r[3] ),
    .A2(_0557_),
    .B(\cnb.data_register_r[4] ),
    .ZN(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1145_ (.A1(_0578_),
    .A2(_0581_),
    .ZN(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1146_ (.A1(_0559_),
    .A2(_0582_),
    .ZN(net34));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1147_ (.I(net34),
    .ZN(net21));
 gf180mcu_fd_sc_mcu7t5v0__buf_20 input10 (.I(a_rst_n),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _1149_ (.A1(_0568_),
    .A2(_0557_),
    .Z(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _1150_ (.A1(\cnb.data_register_r[5] ),
    .A2(\cnb.data_register_r[6] ),
    .A3(_0584_),
    .B(_0559_),
    .ZN(net35));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1151_ (.I(net35),
    .ZN(net22));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _1152_ (.A1(_0252_),
    .A2(_0558_),
    .ZN(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1153_ (.A1(\cnb.data_register_r[5] ),
    .A2(_0574_),
    .B(\cnb.data_register_r[6] ),
    .ZN(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _1154_ (.A1(_0585_),
    .A2(_0586_),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1155_ (.I(net36),
    .ZN(net23));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1156_ (.A1(\cnb.data_register_r[5] ),
    .A2(_0571_),
    .B(\cnb.data_register_r[6] ),
    .ZN(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _1157_ (.A1(_0585_),
    .A2(_0587_),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1158_ (.I(net37),
    .ZN(net24));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1159_ (.A1(_0560_),
    .A2(_0581_),
    .B(_0577_),
    .ZN(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1160_ (.A1(_0559_),
    .A2(_0588_),
    .ZN(net38));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1161_ (.I(net38),
    .ZN(net25));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1162_ (.A1(\cnb.data_register_r[5] ),
    .A2(_0584_),
    .B(\cnb.data_register_r[6] ),
    .ZN(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _1163_ (.A1(_0585_),
    .A2(_0589_),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1164_ (.I(net39),
    .ZN(net26));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1165_ (.A1(\cnb.data_register_r[5] ),
    .A2(_0574_),
    .B(_0559_),
    .C(\cnb.data_register_r[6] ),
    .ZN(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _1166_ (.A1(\cnb.data_register_r[5] ),
    .A2(\cnb.data_register_r[6] ),
    .Z(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _1167_ (.A1(net9),
    .A2(_0568_),
    .A3(net53),
    .A4(_0591_),
    .ZN(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1168_ (.A1(_0590_),
    .A2(_0592_),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1169_ (.I(net40),
    .ZN(net27));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1170_ (.A1(net9),
    .A2(_0571_),
    .B(_0559_),
    .ZN(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _1171_ (.A1(_0585_),
    .A2(_0579_),
    .B1(_0593_),
    .B2(_0560_),
    .ZN(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1172_ (.A1(\cnb.data_register_r[6] ),
    .A2(_0594_),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1173_ (.A1(\cnb.data_register_r[6] ),
    .A2(_0566_),
    .A3(_0567_),
    .ZN(net30));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1174_ (.A1(\cnb.data_register_r[6] ),
    .A2(_0567_),
    .A3(_0573_),
    .ZN(net31));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1175_ (.A1(\cnb.data_register_r[6] ),
    .A2(_0594_),
    .ZN(net41));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1176_ (.A1(_0251_),
    .A2(_0335_),
    .ZN(net43));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1177_ (.A1(_0251_),
    .A2(_0253_),
    .ZN(net44));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1178_ (.A1(_0251_),
    .A2(_0333_),
    .ZN(net45));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1179_ (.A1(_0247_),
    .A2(_0332_),
    .ZN(net104));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _1180_ (.A1(\cnb.data_register_r[9] ),
    .A2(net8),
    .Z(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1181_ (.A1(_0333_),
    .A2(_0595_),
    .ZN(net109));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1182_ (.A1(net104),
    .A2(net109),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1183_ (.A1(_0248_),
    .A2(net8),
    .Z(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1184_ (.I0(_0332_),
    .I1(_0596_),
    .S(\cnb.data_register_r[7] ),
    .Z(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1185_ (.A1(\cnb.data_register_r[8] ),
    .A2(_0597_),
    .ZN(net48));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1186_ (.A1(_0334_),
    .A2(_0248_),
    .ZN(net126));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _1187_ (.A1(net8),
    .A2(net126),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1188_ (.A1(\cnb.data_register_r[8] ),
    .A2(\cnb.data_register_r[9] ),
    .ZN(net67));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1189_ (.A1(net52),
    .A2(net67),
    .ZN(net122));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1190_ (.I(net122),
    .ZN(net113));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _1191_ (.A1(_0252_),
    .A2(net61),
    .A3(net113),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 input9 (.I(a_config_1_in[7]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1193_ (.A1(net8),
    .A2(_0556_),
    .ZN(net50));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _1194_ (.A1(net52),
    .A2(net106),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _1195_ (.A1(net52),
    .A2(net126),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _1196_ (.I(_0333_),
    .ZN(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1197_ (.A1(_0248_),
    .A2(_0599_),
    .Z(net116));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _1198_ (.A1(net8),
    .A2(net116),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1199_ (.I(net64),
    .ZN(net55));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1200_ (.A1(_0453_),
    .A2(_0332_),
    .ZN(net66));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1201_ (.A1(net8),
    .A2(_0599_),
    .B(_0248_),
    .ZN(net56));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _1202_ (.A1(\cnb.data_register_r[9] ),
    .A2(_0453_),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1203_ (.A1(net8),
    .A2(_0333_),
    .B(\cnb.data_register_r[9] ),
    .ZN(net68));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1204_ (.A1(net48),
    .A2(net68),
    .ZN(net58));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1205_ (.I(net61),
    .ZN(net69));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1206_ (.A1(\cnb.data_register_r[9] ),
    .A2(_0333_),
    .Z(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1207_ (.A1(net8),
    .A2(_0600_),
    .ZN(net112));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1208_ (.I(net112),
    .ZN(net121));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1209_ (.A1(_0563_),
    .A2(net121),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_2_0__f_a_clk_dig_in (.I(clknet_0_a_clk_dig_in),
    .Z(clknet_2_0__leaf_a_clk_dig_in));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1211_ (.I(net54),
    .ZN(net63));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1212_ (.I(_0332_),
    .ZN(net65));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1213_ (.A1(net8),
    .A2(_0563_),
    .ZN(net70));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _1214_ (.A1(net52),
    .A2(net116),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _1215_ (.A1(\cnb.data_register_r[7] ),
    .A2(_0558_),
    .Z(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 input8 (.I(a_config_1_in[6]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _1217_ (.A1(_0248_),
    .A2(_0558_),
    .A3(_0599_),
    .B(net52),
    .ZN(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _1218_ (.A1(_0568_),
    .A2(_0603_),
    .Z(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1219_ (.A1(_0591_),
    .A2(_0604_),
    .ZN(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1220_ (.A1(_0601_),
    .A2(_0605_),
    .ZN(net88));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1221_ (.I(net88),
    .ZN(net75));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1222_ (.A1(net9),
    .A2(net121),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1223_ (.A1(_0435_),
    .A2(_0606_),
    .B(_0561_),
    .ZN(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1224_ (.A1(\cnb.data_register_r[4] ),
    .A2(_0607_),
    .B(\cnb.data_register_r[5] ),
    .ZN(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _1225_ (.A1(_0577_),
    .A2(_0585_),
    .Z(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1226_ (.A1(_0608_),
    .A2(_0609_),
    .ZN(net89));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1227_ (.I(net89),
    .ZN(net76));
 gf180mcu_fd_sc_mcu7t5v0__or3_4 _1228_ (.A1(\cnb.data_register_r[3] ),
    .A2(\cnb.data_register_r[4] ),
    .A3(_0603_),
    .Z(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1229_ (.A1(\cnb.data_register_r[3] ),
    .A2(_0603_),
    .B(\cnb.data_register_r[4] ),
    .ZN(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1230_ (.A1(net9),
    .A2(_0611_),
    .ZN(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1231_ (.A1(net9),
    .A2(_0610_),
    .B(_0612_),
    .C(\cnb.data_register_r[5] ),
    .ZN(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1232_ (.A1(_0609_),
    .A2(_0613_),
    .ZN(net90));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1233_ (.I(net90),
    .ZN(net77));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _1234_ (.A1(\cnb.data_register_r[6] ),
    .A2(_0252_),
    .A3(_0604_),
    .B1(_0610_),
    .B2(_0558_),
    .ZN(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1235_ (.A1(_0577_),
    .A2(net9),
    .B1(_0614_),
    .B2(_0560_),
    .ZN(net91));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1236_ (.I(net91),
    .ZN(net78));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _1237_ (.A1(\cnb.data_register_r[3] ),
    .A2(_0603_),
    .Z(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _1238_ (.A1(\cnb.data_register_r[4] ),
    .A2(_0615_),
    .Z(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1239_ (.A1(_0591_),
    .A2(_0616_),
    .ZN(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1240_ (.A1(_0601_),
    .A2(_0617_),
    .ZN(net92));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1241_ (.I(net92),
    .ZN(net79));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1242_ (.A1(\cnb.data_register_r[3] ),
    .A2(_0603_),
    .Z(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _1243_ (.A1(\cnb.data_register_r[4] ),
    .A2(_0618_),
    .Z(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1244_ (.A1(_0591_),
    .A2(_0619_),
    .ZN(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1245_ (.A1(_0601_),
    .A2(_0620_),
    .ZN(net93));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1246_ (.I(net93),
    .ZN(net80));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1247_ (.A1(_0591_),
    .A2(_0610_),
    .ZN(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1248_ (.A1(_0601_),
    .A2(_0621_),
    .ZN(net94));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1249_ (.I(net94),
    .ZN(net81));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1250_ (.A1(\cnb.data_register_r[5] ),
    .A2(_0604_),
    .B(\cnb.data_register_r[6] ),
    .ZN(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1251_ (.A1(_0601_),
    .A2(_0622_),
    .ZN(net95));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1252_ (.I(net95),
    .ZN(net82));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1253_ (.A1(\cnb.data_register_r[5] ),
    .A2(_0616_),
    .B(\cnb.data_register_r[6] ),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1254_ (.A1(_0601_),
    .A2(_0134_),
    .ZN(net96));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1255_ (.I(net96),
    .ZN(net83));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1256_ (.A1(\cnb.data_register_r[5] ),
    .A2(_0619_),
    .B(\cnb.data_register_r[6] ),
    .ZN(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1257_ (.A1(_0601_),
    .A2(_0135_),
    .ZN(net97));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1258_ (.I(net97),
    .ZN(net84));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1259_ (.A1(\cnb.data_register_r[5] ),
    .A2(_0610_),
    .B(\cnb.data_register_r[6] ),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1260_ (.A1(_0601_),
    .A2(_0136_),
    .ZN(net98));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1261_ (.I(net98),
    .ZN(net85));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1262_ (.A1(\cnb.data_register_r[5] ),
    .A2(_0604_),
    .B(_0567_),
    .C(\cnb.data_register_r[6] ),
    .ZN(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _1263_ (.A1(net9),
    .A2(_0449_),
    .A3(net112),
    .Z(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1264_ (.A1(_0137_),
    .A2(_0138_),
    .ZN(net99));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1265_ (.I(net99),
    .ZN(net86));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1266_ (.A1(_0567_),
    .A2(_0612_),
    .ZN(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1267_ (.A1(_0601_),
    .A2(_0611_),
    .B1(_0139_),
    .B2(_0560_),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1268_ (.A1(\cnb.data_register_r[6] ),
    .A2(_0140_),
    .ZN(net87));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _1269_ (.A1(\cnb.data_register_r[6] ),
    .A2(_0140_),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1270_ (.A1(_0253_),
    .A2(_0332_),
    .ZN(net102));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1271_ (.A1(_0332_),
    .A2(_0335_),
    .ZN(net103));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1272_ (.A1(net45),
    .A2(net50),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1273_ (.I0(_0251_),
    .I1(_0595_),
    .S(_0252_),
    .Z(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1274_ (.A1(_0334_),
    .A2(_0141_),
    .ZN(net107));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _1275_ (.A1(net8),
    .A2(net67),
    .Z(net120));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _1276_ (.A1(\cnb.data_register_r[7] ),
    .A2(net54),
    .A3(net120),
    .Z(net108));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1277_ (.A1(_0335_),
    .A2(_0595_),
    .ZN(net110));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1278_ (.I(net8),
    .ZN(net111));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _1279_ (.A1(net8),
    .A2(net57),
    .Z(net123));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1280_ (.I(net123),
    .ZN(net114));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1281_ (.I(_0251_),
    .ZN(net124));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1282_ (.A1(net124),
    .A2(_0563_),
    .ZN(net115));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1283_ (.A1(net8),
    .A2(_0247_),
    .B(_0248_),
    .ZN(net127));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1284_ (.A1(net54),
    .A2(net57),
    .ZN(net117));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1285_ (.I(net120),
    .ZN(net128));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _1286_ (.A1(net52),
    .A2(_0600_),
    .Z(net129));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1287_ (.A1(_0563_),
    .A2(net129),
    .ZN(net118));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_0_a_clk_dig_in (.I(a_clk_dig_in),
    .Z(clknet_0_a_clk_dig_in));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1289_ (.A1(_0251_),
    .A2(_0599_),
    .ZN(net125));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _1290_ (.A1(net52),
    .A2(net57),
    .Z(net130));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1291_ (.A1(\cnb.average_counter_r[0] ),
    .A2(_0373_),
    .ZN(\cnb.next_average_counter_w[0] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1292_ (.A1(_0028_),
    .A2(_0373_),
    .Z(\cnb.next_average_counter_w[1] ));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1293_ (.A1(\cnb.average_counter_r[2] ),
    .A2(_0027_),
    .Z(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1294_ (.A1(_0373_),
    .A2(_0142_),
    .Z(\cnb.next_average_counter_w[2] ));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _1295_ (.A1(\cnb.average_counter_r[2] ),
    .A2(\cnb.average_counter_r[0] ),
    .A3(\cnb.average_counter_r[1] ),
    .Z(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1296_ (.A1(\cnb.average_counter_r[3] ),
    .A2(_0143_),
    .Z(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1297_ (.A1(_0373_),
    .A2(_0144_),
    .Z(\cnb.next_average_counter_w[3] ));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _1298_ (.A1(\cnb.average_counter_r[3] ),
    .A2(\cnb.average_counter_r[2] ),
    .A3(_0027_),
    .Z(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1299_ (.A1(\cnb.average_counter_r[4] ),
    .A2(_0145_),
    .Z(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1300_ (.A1(_0373_),
    .A2(_0146_),
    .Z(\cnb.next_average_counter_w[4] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1301_ (.I0(net1),
    .I1(_0024_),
    .S(_0373_),
    .Z(\cnb.next_average_sum_w[0] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1302_ (.A1(_0026_),
    .A2(_0373_),
    .Z(\cnb.next_average_sum_w[1] ));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1303_ (.A1(\cnb.average_sum_r[2] ),
    .A2(_0025_),
    .Z(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1304_ (.A1(_0373_),
    .A2(_0147_),
    .Z(\cnb.next_average_sum_w[2] ));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _1305_ (.A1(\cnb.average_sum_r[1] ),
    .A2(\cnb.average_sum_r[2] ),
    .A3(_0023_),
    .Z(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1306_ (.A1(\cnb.average_sum_r[3] ),
    .A2(_0148_),
    .Z(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1307_ (.A1(_0373_),
    .A2(_0149_),
    .Z(\cnb.next_average_sum_w[3] ));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _1308_ (.A1(\cnb.average_sum_r[2] ),
    .A2(_0025_),
    .A3(\cnb.average_sum_r[3] ),
    .Z(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1309_ (.A1(\cnb.average_sum_r[4] ),
    .A2(_0150_),
    .Z(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1310_ (.A1(_0373_),
    .A2(_0151_),
    .Z(\cnb.next_average_sum_w[4] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1311_ (.A1(\cnb.is_holding_result_w ),
    .A2(_0347_),
    .Z(\cnb.result_strobe_w ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1312_ (.I(_0503_),
    .ZN(\osr.is_last_sample ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1313_ (.I0(\cnb.result_out[0] ),
    .I1(_0080_),
    .S(_0259_),
    .Z(\osr.next_result_w[0] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1314_ (.I(_0010_),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1315_ (.I0(\cnb.result_out[1] ),
    .I1(_0152_),
    .S(_0259_),
    .Z(\osr.next_result_w[1] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1316_ (.I0(\cnb.result_out[2] ),
    .I1(_0464_),
    .S(_0259_),
    .Z(\osr.next_result_w[2] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1317_ (.A1(\osr.sample_count_r[0] ),
    .A2(_0503_),
    .ZN(\osr.next_sample_count_w[0] ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1318_ (.A1(_0083_),
    .A2(\osr.is_last_sample ),
    .ZN(\osr.next_sample_count_w[1] ));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _1319_ (.A1(_0475_),
    .A2(_0084_),
    .ZN(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1320_ (.A1(_0503_),
    .A2(_0153_),
    .Z(\osr.next_sample_count_w[2] ));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _1321_ (.A1(\osr.sample_count_r[0] ),
    .A2(\osr.sample_count_r[1] ),
    .A3(\osr.sample_count_r[2] ),
    .Z(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1322_ (.A1(\osr.sample_count_r[3] ),
    .A2(_0154_),
    .Z(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1323_ (.A1(_0503_),
    .A2(_0155_),
    .Z(\osr.next_sample_count_w[3] ));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _1324_ (.A1(\osr.sample_count_r[2] ),
    .A2(\osr.sample_count_r[3] ),
    .A3(_0084_),
    .Z(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1325_ (.A1(\osr.sample_count_r[4] ),
    .A2(_0156_),
    .Z(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1326_ (.A1(_0503_),
    .A2(_0157_),
    .Z(\osr.next_sample_count_w[4] ));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _1327_ (.A1(\osr.sample_count_r[0] ),
    .A2(\osr.sample_count_r[1] ),
    .A3(\osr.sample_count_r[2] ),
    .A4(\osr.sample_count_r[3] ),
    .Z(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1328_ (.A1(\osr.sample_count_r[4] ),
    .A2(_0158_),
    .Z(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1329_ (.A1(\osr.sample_count_r[5] ),
    .A2(_0159_),
    .Z(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1330_ (.A1(_0503_),
    .A2(_0160_),
    .Z(\osr.next_sample_count_w[5] ));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _1331_ (.A1(\osr.sample_count_r[4] ),
    .A2(\osr.sample_count_r[5] ),
    .A3(_0156_),
    .Z(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _1332_ (.A1(_0472_),
    .A2(_0161_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1333_ (.A1(_0503_),
    .A2(_0162_),
    .Z(\osr.next_sample_count_w[6] ));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _1334_ (.A1(\osr.sample_count_r[5] ),
    .A2(\osr.sample_count_r[6] ),
    .A3(_0159_),
    .Z(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1335_ (.A1(\osr.sample_count_r[7] ),
    .A2(_0163_),
    .Z(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1336_ (.A1(_0503_),
    .A2(_0164_),
    .Z(\osr.next_sample_count_w[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _1337_ (.A1(\osr.sample_count_r[6] ),
    .A2(\osr.sample_count_r[7] ),
    .A3(_0161_),
    .Z(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _1338_ (.A1(\osr.sample_count_r[8] ),
    .A2(_0165_),
    .Z(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1339_ (.A1(_0503_),
    .A2(_0166_),
    .Z(\osr.next_sample_count_w[8] ));
 gf180mcu_fd_sc_mcu7t5v0__addf_2 _1340_ (.A(net14),
    .B(_0000_),
    .CI(_0001_),
    .CO(_0002_),
    .S(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__addf_2 _1341_ (.A(_0006_),
    .B(_0007_),
    .CI(_0008_),
    .CO(_0009_),
    .S(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _1342_ (.A(_0011_),
    .B(\cnb.average_counter_r[4] ),
    .CO(_0012_),
    .S(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _1343_ (.A(_0014_),
    .B(\cnb.average_counter_r[3] ),
    .CO(_0015_),
    .S(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _1344_ (.A(_0017_),
    .B(\cnb.average_counter_r[2] ),
    .CO(_0018_),
    .S(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _1345_ (.A(_0020_),
    .B(\cnb.average_counter_r[1] ),
    .CO(_0021_),
    .S(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _1346_ (.A(net1),
    .B(\cnb.average_sum_r[0] ),
    .CO(_0023_),
    .S(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _1347_ (.A(\cnb.average_sum_r[1] ),
    .B(_0023_),
    .CO(_0025_),
    .S(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _1348_ (.A(\cnb.average_counter_r[0] ),
    .B(\cnb.average_counter_r[1] ),
    .CO(_0027_),
    .S(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _1349_ (.A(net13),
    .B(net14),
    .CO(_0029_),
    .S(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _1350_ (.A(net72),
    .B(_0031_),
    .CO(_0005_),
    .S(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _1351_ (.A(_0033_),
    .B(_0034_),
    .CO(_0035_),
    .S(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _1352_ (.A(net73),
    .B(_0004_),
    .CO(_0037_),
    .S(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _1353_ (.A(net74),
    .B(_0039_),
    .CO(_0040_),
    .S(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _1354_ (.A(\cnb.data_register_r[3] ),
    .B(_0042_),
    .CO(_0043_),
    .S(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _1355_ (.A(\cnb.data_register_r[4] ),
    .B(_0045_),
    .CO(_0046_),
    .S(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _1356_ (.A(\cnb.data_register_r[5] ),
    .B(_0048_),
    .CO(_0049_),
    .S(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _1357_ (.A(\cnb.data_register_r[6] ),
    .B(_0051_),
    .CO(_0052_),
    .S(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _1358_ (.A(\cnb.data_register_r[7] ),
    .B(_0054_),
    .CO(_0055_),
    .S(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _1359_ (.A(\cnb.data_register_r[6] ),
    .B(_0051_),
    .CO(_0623_),
    .S(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _1360_ (.A(\cnb.data_register_r[8] ),
    .B(_0058_),
    .CO(_0059_),
    .S(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__addh_4 _1361_ (.A(\cnb.result_out[2] ),
    .B(\osr.result_r[2] ),
    .CO(_0061_),
    .S(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _1362_ (.A(\cnb.result_out[1] ),
    .B(\osr.result_r[1] ),
    .CO(_0063_),
    .S(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__addh_4 _1363_ (.A(\cnb.result_out[4] ),
    .B(\osr.result_r[4] ),
    .CO(_0065_),
    .S(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__addh_4 _1364_ (.A(\cnb.result_out[3] ),
    .B(\osr.result_r[3] ),
    .CO(_0067_),
    .S(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _1365_ (.A(\cnb.result_out[6] ),
    .B(\osr.result_r[6] ),
    .CO(_0069_),
    .S(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _1366_ (.A(\cnb.result_out[5] ),
    .B(\osr.result_r[5] ),
    .CO(_0071_),
    .S(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _1367_ (.A(\cnb.result_out[8] ),
    .B(\osr.result_r[8] ),
    .CO(_0073_),
    .S(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _1368_ (.A(\cnb.result_out[7] ),
    .B(\osr.result_r[7] ),
    .CO(_0075_),
    .S(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _1369_ (.A(\cnb.result_out[9] ),
    .B(\osr.result_r[9] ),
    .CO(_0077_),
    .S(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _1370_ (.A(\cnb.result_out[0] ),
    .B(\osr.result_r[0] ),
    .CO(_0079_),
    .S(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _1371_ (.A(\osr.sample_count_r[0] ),
    .B(_0081_),
    .CO(_0082_),
    .S(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__addh_2 _1372_ (.A(\osr.sample_count_r[0] ),
    .B(\osr.sample_count_r[1] ),
    .CO(_0084_),
    .S(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__tieh _1375__4 (.Z(a_nmatrix_c0_out_n));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input7 (.I(a_config_1_in[5]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input6 (.I(a_config_1_in[4]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input5 (.I(a_config_1_in[3]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input4 (.I(a_config_1_in[2]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input3 (.I(a_config_1_in[1]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input2 (.I(a_config_1_in[0]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input1 (.I(a_comparator_in),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_2_3__f_a_clk_dig_in (.I(clknet_0_a_clk_dig_in),
    .Z(clknet_2_3__leaf_a_clk_dig_in));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_2_1__f_a_clk_dig_in (.I(clknet_0_a_clk_dig_in),
    .Z(clknet_2_1__leaf_a_clk_dig_in));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_2_2__f_a_clk_dig_in (.I(clknet_0_a_clk_dig_in),
    .Z(clknet_2_2__leaf_a_clk_dig_in));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_4 \cnb.average_counter_r[0]$_DFF_PN1_  (.D(\cnb.next_average_counter_w[0] ),
    .SETN(net10),
    .CLK(clknet_2_0__leaf_a_clk_dig_in),
    .Q(\cnb.average_counter_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.average_counter_r[1]$_DFF_PN0_  (.D(\cnb.next_average_counter_w[1] ),
    .RN(net10),
    .CLK(clknet_2_0__leaf_a_clk_dig_in),
    .Q(\cnb.average_counter_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.average_counter_r[2]$_DFF_PN0_  (.D(\cnb.next_average_counter_w[2] ),
    .RN(net10),
    .CLK(clknet_2_0__leaf_a_clk_dig_in),
    .Q(\cnb.average_counter_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.average_counter_r[3]$_DFF_PN0_  (.D(\cnb.next_average_counter_w[3] ),
    .RN(net10),
    .CLK(clknet_2_1__leaf_a_clk_dig_in),
    .Q(\cnb.average_counter_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.average_counter_r[4]$_DFF_PN0_  (.D(\cnb.next_average_counter_w[4] ),
    .RN(net10),
    .CLK(clknet_2_0__leaf_a_clk_dig_in),
    .Q(\cnb.average_counter_r[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.average_sum_r[0]$_DFF_PN0_  (.D(\cnb.next_average_sum_w[0] ),
    .RN(net10),
    .CLK(clknet_2_0__leaf_a_clk_dig_in),
    .Q(\cnb.average_sum_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.average_sum_r[1]$_DFF_PN0_  (.D(\cnb.next_average_sum_w[1] ),
    .RN(net10),
    .CLK(clknet_2_0__leaf_a_clk_dig_in),
    .Q(\cnb.average_sum_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.average_sum_r[2]$_DFF_PN0_  (.D(\cnb.next_average_sum_w[2] ),
    .RN(net10),
    .CLK(clknet_2_0__leaf_a_clk_dig_in),
    .Q(\cnb.average_sum_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.average_sum_r[3]$_DFF_PN0_  (.D(\cnb.next_average_sum_w[3] ),
    .RN(net10),
    .CLK(clknet_2_0__leaf_a_clk_dig_in),
    .Q(\cnb.average_sum_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.average_sum_r[4]$_DFF_PN0_  (.D(\cnb.next_average_sum_w[4] ),
    .RN(net10),
    .CLK(clknet_2_0__leaf_a_clk_dig_in),
    .Q(\cnb.average_sum_r[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.conv_finished_r$_DFF_PN0_  (.D(\cnb.result_strobe_w ),
    .RN(net10),
    .CLK(clknet_2_0__leaf_a_clk_dig_in),
    .Q(\cnb.conv_finished_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.data_register_r[0]$_DFFE_PN0P_  (.D(_0085_),
    .RN(net10),
    .CLK(clknet_2_1__leaf_a_clk_dig_in),
    .Q(net72));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.data_register_r[1]$_DFFE_PN0P_  (.D(_0086_),
    .RN(net10),
    .CLK(clknet_2_1__leaf_a_clk_dig_in),
    .Q(net73));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.data_register_r[2]$_DFFE_PN0P_  (.D(_0087_),
    .RN(net10),
    .CLK(clknet_2_3__leaf_a_clk_dig_in),
    .Q(net74));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.data_register_r[3]$_DFFE_PN0P_  (.D(_0088_),
    .RN(net10),
    .CLK(clknet_2_3__leaf_a_clk_dig_in),
    .Q(\cnb.data_register_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.data_register_r[4]$_DFFE_PN0P_  (.D(_0089_),
    .RN(net10),
    .CLK(clknet_2_3__leaf_a_clk_dig_in),
    .Q(\cnb.data_register_r[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.data_register_r[5]$_DFFE_PN0P_  (.D(_0090_),
    .RN(net10),
    .CLK(clknet_2_3__leaf_a_clk_dig_in),
    .Q(\cnb.data_register_r[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.data_register_r[6]$_DFFE_PN0P_  (.D(_0091_),
    .RN(net10),
    .CLK(clknet_2_3__leaf_a_clk_dig_in),
    .Q(\cnb.data_register_r[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.data_register_r[7]$_DFFE_PN0P_  (.D(_0092_),
    .RN(net10),
    .CLK(clknet_2_3__leaf_a_clk_dig_in),
    .Q(\cnb.data_register_r[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.data_register_r[8]$_DFFE_PN0P_  (.D(_0093_),
    .RN(net10),
    .CLK(clknet_2_3__leaf_a_clk_dig_in),
    .Q(\cnb.data_register_r[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_4 \cnb.data_register_r[9]$_DFFE_PN1P_  (.D(_0094_),
    .SETN(net10),
    .CLK(clknet_2_2__leaf_a_clk_dig_in),
    .Q(\cnb.data_register_r[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.result_out[0]$_DFFE_PN0P_  (.D(_0095_),
    .RN(net10),
    .CLK(clknet_2_1__leaf_a_clk_dig_in),
    .Q(\cnb.result_out[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.result_out[1]$_DFFE_PN0P_  (.D(_0096_),
    .RN(net10),
    .CLK(clknet_2_1__leaf_a_clk_dig_in),
    .Q(\cnb.result_out[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.result_out[2]$_DFFE_PN0P_  (.D(_0097_),
    .RN(net10),
    .CLK(clknet_2_1__leaf_a_clk_dig_in),
    .Q(\cnb.result_out[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.result_out[3]$_DFFE_PN0P_  (.D(_0098_),
    .RN(net10),
    .CLK(clknet_2_1__leaf_a_clk_dig_in),
    .Q(\cnb.result_out[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.result_out[4]$_DFFE_PN0P_  (.D(_0099_),
    .RN(net10),
    .CLK(clknet_2_1__leaf_a_clk_dig_in),
    .Q(\cnb.result_out[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.result_out[5]$_DFFE_PN0P_  (.D(_0100_),
    .RN(net10),
    .CLK(clknet_2_3__leaf_a_clk_dig_in),
    .Q(\cnb.result_out[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.result_out[6]$_DFFE_PN0P_  (.D(_0101_),
    .RN(net10),
    .CLK(clknet_2_1__leaf_a_clk_dig_in),
    .Q(\cnb.result_out[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.result_out[7]$_DFFE_PN0P_  (.D(_0102_),
    .RN(net10),
    .CLK(clknet_2_1__leaf_a_clk_dig_in),
    .Q(\cnb.result_out[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.result_out[8]$_DFFE_PN0P_  (.D(_0103_),
    .RN(net10),
    .CLK(clknet_2_3__leaf_a_clk_dig_in),
    .Q(\cnb.result_out[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.result_out[9]$_DFFE_PN0P_  (.D(_0104_),
    .RN(net10),
    .CLK(clknet_2_1__leaf_a_clk_dig_in),
    .Q(\cnb.result_out[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.sampled_avg_control_r[0]$_DFFE_PN0P_  (.D(_0105_),
    .RN(net10),
    .CLK(clknet_2_0__leaf_a_clk_dig_in),
    .Q(\cnb.sampled_avg_control_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.sampled_avg_control_r[1]$_DFFE_PN0P_  (.D(_0106_),
    .RN(net10),
    .CLK(clknet_2_0__leaf_a_clk_dig_in),
    .Q(\cnb.sampled_avg_control_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.sampled_avg_control_r[2]$_DFFE_PN0P_  (.D(_0107_),
    .RN(net10),
    .CLK(clknet_2_0__leaf_a_clk_dig_in),
    .Q(\cnb.sampled_avg_control_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_4 \cnb.shift_register_r[0]$_DFFE_PN1N_  (.D(_0108_),
    .SETN(net10),
    .CLK(clknet_2_0__leaf_a_clk_dig_in),
    .Q(net139));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.shift_register_r[10]$_DFFE_PN0N_  (.D(_0109_),
    .RN(net10),
    .CLK(clknet_2_2__leaf_a_clk_dig_in),
    .Q(\cnb.shift_register_r[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.shift_register_r[11]$_DFFE_PN0N_  (.D(_0110_),
    .RN(net10),
    .CLK(clknet_2_2__leaf_a_clk_dig_in),
    .Q(\cnb.shift_register_r[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.shift_register_r[12]$_DFFE_PN0N_  (.D(_0111_),
    .RN(net10),
    .CLK(clknet_2_2__leaf_a_clk_dig_in),
    .Q(\cnb.shift_register_r[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.shift_register_r[13]$_DFFE_PN0N_  (.D(_0112_),
    .RN(net10),
    .CLK(clknet_2_2__leaf_a_clk_dig_in),
    .Q(\cnb.shift_register_r[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.shift_register_r[14]$_DFFE_PN0N_  (.D(_0113_),
    .RN(net10),
    .CLK(clknet_2_2__leaf_a_clk_dig_in),
    .Q(\cnb.shift_register_r[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.shift_register_r[1]$_DFFE_PN0N_  (.D(_0114_),
    .RN(net10),
    .CLK(clknet_2_0__leaf_a_clk_dig_in),
    .Q(\cnb.is_holding_result_w ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.shift_register_r[2]$_DFFE_PN0N_  (.D(_0115_),
    .RN(net10),
    .CLK(clknet_2_1__leaf_a_clk_dig_in),
    .Q(\cnb.shift_register_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.shift_register_r[3]$_DFFE_PN0N_  (.D(_0116_),
    .RN(net10),
    .CLK(clknet_2_0__leaf_a_clk_dig_in),
    .Q(\cnb.shift_register_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.shift_register_r[4]$_DFFE_PN0N_  (.D(_0117_),
    .RN(net10),
    .CLK(clknet_2_2__leaf_a_clk_dig_in),
    .Q(\cnb.shift_register_r[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.shift_register_r[5]$_DFFE_PN0N_  (.D(_0118_),
    .RN(net10),
    .CLK(clknet_2_2__leaf_a_clk_dig_in),
    .Q(\cnb.shift_register_r[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.shift_register_r[6]$_DFFE_PN0N_  (.D(_0119_),
    .RN(net10),
    .CLK(clknet_2_2__leaf_a_clk_dig_in),
    .Q(\cnb.shift_register_r[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.shift_register_r[7]$_DFFE_PN0N_  (.D(_0120_),
    .RN(net10),
    .CLK(clknet_2_2__leaf_a_clk_dig_in),
    .Q(\cnb.shift_register_r[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.shift_register_r[8]$_DFFE_PN0N_  (.D(_0121_),
    .RN(net10),
    .CLK(clknet_2_2__leaf_a_clk_dig_in),
    .Q(\cnb.shift_register_r[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \cnb.shift_register_r[9]$_DFFE_PN0N_  (.D(_0122_),
    .RN(net10),
    .CLK(clknet_2_2__leaf_a_clk_dig_in),
    .Q(\cnb.shift_register_r[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \osr.data_valid_r$_DFF_PN0_  (.D(\osr.is_last_sample ),
    .RN(net10),
    .CLK(\cnb.conv_finished_r ),
    .Q(\osr.data_valid_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \osr.osr_mode_r[0]$_DFFE_PN0P_  (.D(_0123_),
    .RN(net10),
    .CLK(\cnb.conv_finished_r ),
    .Q(\osr.osr_mode_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \osr.osr_mode_r[1]$_DFFE_PN0P_  (.D(_0124_),
    .RN(net10),
    .CLK(\cnb.conv_finished_r ),
    .Q(\osr.osr_mode_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \osr.osr_mode_r[2]$_DFFE_PN0P_  (.D(_0125_),
    .RN(net10),
    .CLK(\cnb.conv_finished_r ),
    .Q(\osr.osr_mode_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \osr.output_r[2]$_DFFE_PN0P_  (.D(_0126_),
    .RN(net10),
    .CLK(\cnb.conv_finished_r ),
    .Q(net131));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \osr.output_r[3]$_DFFE_PN0P_  (.D(_0127_),
    .RN(net10),
    .CLK(\cnb.conv_finished_r ),
    .Q(net132));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \osr.output_r[4]$_DFFE_PN0P_  (.D(_0128_),
    .RN(net10),
    .CLK(\cnb.conv_finished_r ),
    .Q(net133));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \osr.output_r[5]$_DFFE_PN0P_  (.D(_0129_),
    .RN(net10),
    .CLK(\cnb.conv_finished_r ),
    .Q(net134));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \osr.output_r[6]$_DFFE_PN0P_  (.D(_0130_),
    .RN(net10),
    .CLK(\cnb.conv_finished_r ),
    .Q(net135));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \osr.output_r[7]$_DFFE_PN0P_  (.D(_0131_),
    .RN(net10),
    .CLK(\cnb.conv_finished_r ),
    .Q(net136));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \osr.output_r[8]$_DFFE_PN0P_  (.D(_0132_),
    .RN(net10),
    .CLK(\cnb.conv_finished_r ),
    .Q(net137));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \osr.output_r[9]$_DFFE_PN0P_  (.D(_0133_),
    .RN(net10),
    .CLK(\cnb.conv_finished_r ),
    .Q(net138));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \osr.result_r[0]$_DFF_PN0_  (.D(\osr.next_result_w[0] ),
    .RN(net10),
    .CLK(\cnb.conv_finished_r ),
    .Q(\osr.result_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \osr.result_r[10]$_DFF_PN0_  (.D(\osr.next_result_w[10] ),
    .RN(net10),
    .CLK(\cnb.conv_finished_r ),
    .Q(\osr.result_r[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \osr.result_r[11]$_DFF_PN0_  (.D(\osr.next_result_w[11] ),
    .RN(net10),
    .CLK(\cnb.conv_finished_r ),
    .Q(\osr.result_r[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \osr.result_r[12]$_DFF_PN0_  (.D(\osr.next_result_w[12] ),
    .RN(net10),
    .CLK(\cnb.conv_finished_r ),
    .Q(\osr.result_r[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \osr.result_r[13]$_DFF_PN0_  (.D(\osr.next_result_w[13] ),
    .RN(net10),
    .CLK(\cnb.conv_finished_r ),
    .Q(\osr.result_r[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \osr.result_r[14]$_DFF_PN0_  (.D(\osr.next_result_w[14] ),
    .RN(net10),
    .CLK(\cnb.conv_finished_r ),
    .Q(\osr.result_r[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \osr.result_r[15]$_DFF_PN0_  (.D(\osr.next_result_w[15] ),
    .RN(net10),
    .CLK(\cnb.conv_finished_r ),
    .Q(\osr.result_r[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \osr.result_r[1]$_DFF_PN0_  (.D(\osr.next_result_w[1] ),
    .RN(net10),
    .CLK(\cnb.conv_finished_r ),
    .Q(\osr.result_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \osr.result_r[2]$_DFF_PN0_  (.D(\osr.next_result_w[2] ),
    .RN(net10),
    .CLK(\cnb.conv_finished_r ),
    .Q(\osr.result_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \osr.result_r[3]$_DFF_PN0_  (.D(\osr.next_result_w[3] ),
    .RN(net10),
    .CLK(\cnb.conv_finished_r ),
    .Q(\osr.result_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \osr.result_r[4]$_DFF_PN0_  (.D(\osr.next_result_w[4] ),
    .RN(net10),
    .CLK(\cnb.conv_finished_r ),
    .Q(\osr.result_r[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \osr.result_r[5]$_DFF_PN0_  (.D(\osr.next_result_w[5] ),
    .RN(net10),
    .CLK(\cnb.conv_finished_r ),
    .Q(\osr.result_r[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \osr.result_r[6]$_DFF_PN0_  (.D(\osr.next_result_w[6] ),
    .RN(net10),
    .CLK(\cnb.conv_finished_r ),
    .Q(\osr.result_r[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \osr.result_r[7]$_DFF_PN0_  (.D(\osr.next_result_w[7] ),
    .RN(net10),
    .CLK(\cnb.conv_finished_r ),
    .Q(\osr.result_r[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \osr.result_r[8]$_DFF_PN0_  (.D(\osr.next_result_w[8] ),
    .RN(net10),
    .CLK(\cnb.conv_finished_r ),
    .Q(\osr.result_r[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \osr.result_r[9]$_DFF_PN0_  (.D(\osr.next_result_w[9] ),
    .RN(net10),
    .CLK(\cnb.conv_finished_r ),
    .Q(\osr.result_r[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_4 \osr.sample_count_r[0]$_DFF_PN1_  (.D(\osr.next_sample_count_w[0] ),
    .SETN(net10),
    .CLK(\cnb.conv_finished_r ),
    .Q(\osr.sample_count_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \osr.sample_count_r[1]$_DFF_PN0_  (.D(\osr.next_sample_count_w[1] ),
    .RN(net10),
    .CLK(\cnb.conv_finished_r ),
    .Q(\osr.sample_count_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \osr.sample_count_r[2]$_DFF_PN0_  (.D(\osr.next_sample_count_w[2] ),
    .RN(net10),
    .CLK(\cnb.conv_finished_r ),
    .Q(\osr.sample_count_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \osr.sample_count_r[3]$_DFF_PN0_  (.D(\osr.next_sample_count_w[3] ),
    .RN(net10),
    .CLK(\cnb.conv_finished_r ),
    .Q(\osr.sample_count_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \osr.sample_count_r[4]$_DFF_PN0_  (.D(\osr.next_sample_count_w[4] ),
    .RN(net10),
    .CLK(\cnb.conv_finished_r ),
    .Q(\osr.sample_count_r[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \osr.sample_count_r[5]$_DFF_PN0_  (.D(\osr.next_sample_count_w[5] ),
    .RN(net10),
    .CLK(\cnb.conv_finished_r ),
    .Q(\osr.sample_count_r[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \osr.sample_count_r[6]$_DFF_PN0_  (.D(\osr.next_sample_count_w[6] ),
    .RN(net10),
    .CLK(\cnb.conv_finished_r ),
    .Q(\osr.sample_count_r[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \osr.sample_count_r[7]$_DFF_PN0_  (.D(\osr.next_sample_count_w[7] ),
    .RN(net10),
    .CLK(\cnb.conv_finished_r ),
    .Q(\osr.sample_count_r[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \osr.sample_count_r[8]$_DFF_PN0_  (.D(\osr.next_sample_count_w[8] ),
    .RN(net10),
    .CLK(\cnb.conv_finished_r ),
    .Q(\osr.sample_count_r[8] ));
 gf180mcu_fd_sc_mcu7t5v0__tiel _1379__1 (.ZN(a_pmatrix_c0_out_n));
 gf180mcu_fd_sc_mcu7t5v0__tiel _1380__2 (.ZN(a_result_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _1381__3 (.ZN(a_result_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Left_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Left_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Left_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Left_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Left_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Left_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Left_109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_166 ();
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output30 (.I(net30),
    .Z(a_nmatrix_col_out_n[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output31 (.I(net31),
    .Z(a_nmatrix_col_out_n[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output32 (.I(net32),
    .Z(a_nmatrix_col_out_n[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output33 (.I(net33),
    .Z(a_nmatrix_col_out_n[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output34 (.I(net34),
    .Z(a_nmatrix_col_out_n[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output35 (.I(net35),
    .Z(a_nmatrix_col_out_n[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output36 (.I(net36),
    .Z(a_nmatrix_col_out_n[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output37 (.I(net37),
    .Z(a_nmatrix_col_out_n[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output38 (.I(net38),
    .Z(a_nmatrix_col_out_n[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output39 (.I(net39),
    .Z(a_nmatrix_col_out_n[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output40 (.I(net40),
    .Z(a_nmatrix_col_out_n[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output41 (.I(net41),
    .Z(a_nmatrix_col_out_n[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output42 (.I(net42),
    .Z(a_nmatrix_row_out_n[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output43 (.I(net43),
    .Z(a_nmatrix_row_out_n[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output44 (.I(net44),
    .Z(a_nmatrix_row_out_n[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output45 (.I(net45),
    .Z(a_nmatrix_row_out_n[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output46 (.I(net46),
    .Z(a_nmatrix_row_out_n[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output47 (.I(net47),
    .Z(a_nmatrix_row_out_n[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output48 (.I(net48),
    .Z(a_nmatrix_row_out_n[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output49 (.I(net49),
    .Z(a_nmatrix_row_out_n[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output50 (.I(net50),
    .Z(a_nmatrix_row_out_n[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output51 (.I(net51),
    .Z(a_nmatrix_row_out_n[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output52 (.I(net52),
    .Z(a_nmatrix_rowoff_out_n[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output53 (.I(net53),
    .Z(a_nmatrix_rowoff_out_n[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output54 (.I(net54),
    .Z(a_nmatrix_rowoff_out_n[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output55 (.I(net55),
    .Z(a_nmatrix_rowoff_out_n[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output56 (.I(net56),
    .Z(a_nmatrix_rowoff_out_n[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output57 (.I(net57),
    .Z(a_nmatrix_rowoff_out_n[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output58 (.I(net58),
    .Z(a_nmatrix_rowoff_out_n[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output59 (.I(net59),
    .Z(a_nmatrix_rowoff_out_n[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output60 (.I(net8),
    .Z(a_nmatrix_rowoff_out_n[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output61 (.I(net61),
    .Z(a_nmatrix_rowoff_out_n[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output62 (.I(net62),
    .Z(a_nmatrix_rowon_out_n[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output63 (.I(net63),
    .Z(a_nmatrix_rowon_out_n[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output64 (.I(net64),
    .Z(a_nmatrix_rowon_out_n[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output65 (.I(net65),
    .Z(a_nmatrix_rowon_out_n[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output66 (.I(net66),
    .Z(a_nmatrix_rowon_out_n[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output67 (.I(net67),
    .Z(a_nmatrix_rowon_out_n[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output68 (.I(net68),
    .Z(a_nmatrix_rowon_out_n[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output69 (.I(net69),
    .Z(a_nmatrix_rowon_out_n[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output70 (.I(net70),
    .Z(a_nmatrix_rowon_out_n[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output71 (.I(net71),
    .Z(a_nmatrix_rowon_out_n[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output72 (.I(net72),
    .Z(a_pmatrix_bincap_out_n[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output73 (.I(net73),
    .Z(a_pmatrix_bincap_out_n[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output74 (.I(net74),
    .Z(a_pmatrix_bincap_out_n[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output75 (.I(net75),
    .Z(a_pmatrix_col_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output76 (.I(net76),
    .Z(a_pmatrix_col_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output77 (.I(net77),
    .Z(a_pmatrix_col_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output78 (.I(net78),
    .Z(a_pmatrix_col_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output79 (.I(net79),
    .Z(a_pmatrix_col_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output80 (.I(net80),
    .Z(a_pmatrix_col_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output81 (.I(net81),
    .Z(a_pmatrix_col_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output82 (.I(net82),
    .Z(a_pmatrix_col_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output83 (.I(net83),
    .Z(a_pmatrix_col_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output84 (.I(net84),
    .Z(a_pmatrix_col_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output85 (.I(net85),
    .Z(a_pmatrix_col_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output86 (.I(net86),
    .Z(a_pmatrix_col_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output87 (.I(net87),
    .Z(a_pmatrix_col_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output88 (.I(net88),
    .Z(a_pmatrix_col_out_n[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output89 (.I(net89),
    .Z(a_pmatrix_col_out_n[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output90 (.I(net90),
    .Z(a_pmatrix_col_out_n[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output91 (.I(net91),
    .Z(a_pmatrix_col_out_n[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output92 (.I(net92),
    .Z(a_pmatrix_col_out_n[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output93 (.I(net93),
    .Z(a_pmatrix_col_out_n[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output94 (.I(net94),
    .Z(a_pmatrix_col_out_n[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output95 (.I(net95),
    .Z(a_pmatrix_col_out_n[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output96 (.I(net96),
    .Z(a_pmatrix_col_out_n[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output97 (.I(net97),
    .Z(a_pmatrix_col_out_n[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output98 (.I(net98),
    .Z(a_pmatrix_col_out_n[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output99 (.I(net99),
    .Z(a_pmatrix_col_out_n[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output100 (.I(net100),
    .Z(a_pmatrix_col_out_n[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output101 (.I(net101),
    .Z(a_pmatrix_row_out_n[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output102 (.I(net102),
    .Z(a_pmatrix_row_out_n[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output103 (.I(net103),
    .Z(a_pmatrix_row_out_n[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output104 (.I(net104),
    .Z(a_pmatrix_row_out_n[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output105 (.I(net105),
    .Z(a_pmatrix_row_out_n[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output106 (.I(net106),
    .Z(a_pmatrix_row_out_n[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output107 (.I(net107),
    .Z(a_pmatrix_row_out_n[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output108 (.I(net108),
    .Z(a_pmatrix_row_out_n[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output109 (.I(net109),
    .Z(a_pmatrix_row_out_n[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output110 (.I(net110),
    .Z(a_pmatrix_row_out_n[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output111 (.I(net111),
    .Z(a_pmatrix_rowoff_out_n[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output112 (.I(net112),
    .Z(a_pmatrix_rowoff_out_n[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output113 (.I(net113),
    .Z(a_pmatrix_rowoff_out_n[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output114 (.I(net114),
    .Z(a_pmatrix_rowoff_out_n[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output115 (.I(net115),
    .Z(a_pmatrix_rowoff_out_n[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output116 (.I(net116),
    .Z(a_pmatrix_rowoff_out_n[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output117 (.I(net117),
    .Z(a_pmatrix_rowoff_out_n[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output118 (.I(net118),
    .Z(a_pmatrix_rowoff_out_n[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output119 (.I(net8),
    .Z(a_pmatrix_rowoff_out_n[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output120 (.I(net120),
    .Z(a_pmatrix_rowoff_out_n[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output121 (.I(net121),
    .Z(a_pmatrix_rowon_out_n[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output122 (.I(net122),
    .Z(a_pmatrix_rowon_out_n[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output123 (.I(net123),
    .Z(a_pmatrix_rowon_out_n[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output124 (.I(net124),
    .Z(a_pmatrix_rowon_out_n[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output125 (.I(net125),
    .Z(a_pmatrix_rowon_out_n[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output126 (.I(net126),
    .Z(a_pmatrix_rowon_out_n[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output127 (.I(net127),
    .Z(a_pmatrix_rowon_out_n[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output128 (.I(net128),
    .Z(a_pmatrix_rowon_out_n[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output129 (.I(net129),
    .Z(a_pmatrix_rowon_out_n[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output130 (.I(net130),
    .Z(a_pmatrix_rowon_out_n[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output131 (.I(net131),
    .Z(a_result_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output132 (.I(net132),
    .Z(a_result_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output133 (.I(net133),
    .Z(a_result_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output134 (.I(net134),
    .Z(a_result_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output135 (.I(net135),
    .Z(a_result_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output136 (.I(net136),
    .Z(a_result_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output137 (.I(net137),
    .Z(a_result_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output138 (.I(net138),
    .Z(a_result_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output139 (.I(net139),
    .Z(a_sample_matrix_out));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output140 (.I(net12),
    .Z(a_sample_matrix_out_n));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output141 (.I(net139),
    .Z(a_sample_switch_out));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 output142 (.I(net12),
    .Z(a_sample_switch_out_n));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 clkload0 (.I(clknet_2_1__leaf_a_clk_dig_in));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 clkload1 (.I(clknet_2_2__leaf_a_clk_dig_in));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkload2 (.I(clknet_2_3__leaf_a_clk_dig_in));
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_0_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_0_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_0_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_0_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_0_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_0_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_0_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_0_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_0_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_0_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_1_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_1_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_1_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_1_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_1_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_1_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_1_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_1_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_1_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_1_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_1_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_2_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_2_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_2_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_2_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_2_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_2_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_3_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_3_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_3_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_3_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_3_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_3_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_3_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_3_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_4_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_4_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_4_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_4_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_4_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_4_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_5_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_5_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_5_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_5_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_5_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_5_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_5_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_5_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_6_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_6_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_6_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_6_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_6_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_6_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_6_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_6_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_6_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_6_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_6_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_7_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_7_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_7_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_7_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_7_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_7_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_7_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_7_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_7_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_7_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_7_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_7_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_7_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_7_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_8_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_8_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_8_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_8_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_8_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_8_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_8_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_8_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_8_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_8_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_9_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_9_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_9_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_9_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_9_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_9_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_9_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_9_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_9_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_9_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_10_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_10_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_10_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_10_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_10_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_10_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_10_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_10_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_10_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_10_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_11_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_11_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_11_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_11_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_11_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_11_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_11_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_11_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_11_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_11_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_11_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_11_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_11_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_11_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_12_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_12_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_12_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_12_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_12_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_12_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_12_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_12_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_12_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_13_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_13_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_13_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_13_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_13_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_13_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_13_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_13_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_13_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_14_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_14_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_14_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_14_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_14_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_15_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_15_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_15_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_15_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_15_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_15_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_15_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_15_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_15_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_15_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_15_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_16_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_16_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_16_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_16_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_16_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_16_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_16_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_16_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_16_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_16_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_17_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_17_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_17_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_17_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_17_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_17_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_17_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_17_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_18_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_18_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_18_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_18_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_18_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_18_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_18_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_18_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_18_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_19_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_19_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_19_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_19_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_19_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_19_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_19_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_19_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_19_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_19_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_19_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_19_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_20_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_20_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_20_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_20_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_20_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_20_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_20_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_20_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_21_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_21_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_21_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_21_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_21_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_21_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_22_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_22_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_22_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_22_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_23_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_23_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_23_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_23_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_23_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_23_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_23_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_23_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_23_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_23_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_23_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_23_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_23_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_24_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_24_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_24_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_24_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_24_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_24_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_24_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_24_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_24_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_24_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_24_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_24_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_24_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_24_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_24_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_24_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_25_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_25_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_25_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_25_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_25_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_25_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_25_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_26_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_26_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_26_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_26_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_26_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_26_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_26_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_26_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_26_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_27_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_27_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_27_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_27_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_27_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_27_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_27_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_27_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_27_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_28_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_28_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_28_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_28_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_28_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_28_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_28_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_28_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_28_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_28_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_28_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_28_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_28_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_28_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_28_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_29_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_29_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_29_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_29_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_29_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_29_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_29_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_29_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_29_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_29_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_29_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_29_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_30_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_30_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_30_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_30_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_30_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_30_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_30_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_31_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_31_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_31_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_31_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_31_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_31_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_31_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_31_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_31_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_31_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_31_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_31_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_31_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_31_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_32_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_32_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_32_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_32_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_32_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_32_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_32_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_33_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_33_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_33_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_33_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_33_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_33_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_33_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_33_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_33_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_34_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_34_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_34_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_34_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_34_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_34_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_34_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_34_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_34_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_34_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_34_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_34_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_34_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_34_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_34_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_34_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_35_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_35_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_35_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_35_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_35_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_36_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_36_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_36_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_36_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_36_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_36_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_37_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_37_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_37_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_37_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_37_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_37_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_38_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_38_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_38_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_38_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_38_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_38_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_38_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_39_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_39_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_39_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_39_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_39_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_39_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_39_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_39_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_39_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_39_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_39_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_40_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_40_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_40_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_40_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_40_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_40_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_40_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_40_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_40_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_41_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_41_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_41_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_41_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_41_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_41_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_41_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_41_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_41_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_41_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_41_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_41_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_41_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_42_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_42_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_42_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_42_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_42_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_42_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_42_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_42_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_42_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_43_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_43_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_43_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_43_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_43_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_43_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_43_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_43_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_43_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_44_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_44_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_44_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_44_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_44_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_44_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_44_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_44_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_44_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_45_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_45_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_45_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_45_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_45_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_45_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_45_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_45_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_46_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_46_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_46_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_46_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_46_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_46_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_46_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_46_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_46_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_46_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_47_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_47_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_47_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_47_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_47_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_47_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_47_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_47_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_47_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_47_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_47_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_48_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_48_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_48_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_48_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_48_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_48_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_48_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_48_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_48_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_48_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_48_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_49_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_49_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_49_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_49_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_49_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_49_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_49_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_49_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_49_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_49_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_49_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_49_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_49_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_50_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_50_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_50_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_50_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_50_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_50_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_50_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_50_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_50_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_50_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_51_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_51_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_51_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_51_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_51_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_51_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_51_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_51_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_51_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_51_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_51_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_52_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_52_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_52_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_52_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_52_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_52_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_52_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_52_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_52_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_52_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_53_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_53_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_53_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_53_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_53_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_53_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_53_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_53_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_53_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_53_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_53_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_64 FILLER_54_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_32 FILLER_54_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_54_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_54_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_8 FILLER_54_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_54_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_16 FILLER_54_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_4 FILLER_54_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_391 ();
endmodule
