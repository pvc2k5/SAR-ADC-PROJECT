module adc_clkgen_with_edgedetect (VDD,
    VSS,
    clk_comp_out,
    clk_dig_out,
    ena_in,
    enable_dlycontrol_in,
    ndecision_finish_in,
    sample_n_in,
    sample_n_out,
    sample_p_in,
    sample_p_out,
    start_conv_in,
    dlycontrol1_in,
    dlycontrol2_in,
    dlycontrol3_in,
    dlycontrol4_in);
 input VDD;
 input VSS;
 output clk_comp_out;
 output clk_dig_out;
 input ena_in;
 input enable_dlycontrol_in;
 input ndecision_finish_in;
 input sample_n_in;
 output sample_n_out;
 input sample_p_in;
 output sample_p_out;
 input start_conv_in;
 input [4:0] dlycontrol1_in;
 input [4:0] dlycontrol2_in;
 input [4:0] dlycontrol3_in;
 input [5:0] dlycontrol4_in;

 wire \clkgen.clk_comp_out ;
 wire \clkgen.clk_dig_delayed_w ;
 wire \clkgen.clk_dig_out ;
 wire \clkgen.delay_155ns_1.bypass_enable_w[0] ;
 wire \clkgen.delay_155ns_1.bypass_enable_w[1] ;
 wire \clkgen.delay_155ns_1.bypass_enable_w[2] ;
 wire \clkgen.delay_155ns_1.bypass_enable_w[3] ;
 wire \clkgen.delay_155ns_1.bypass_enable_w[4] ;
 wire \clkgen.delay_155ns_1.enable_dlycontrol_w ;
 wire \clkgen.delay_155ns_1.genblk1[0].dly_binary.bypass_in ;
 wire \clkgen.delay_155ns_1.genblk1[0].dly_binary.in ;
 wire \clkgen.delay_155ns_1.genblk1[0].dly_binary.out ;
 wire \clkgen.delay_155ns_1.genblk1[0].dly_binary.signal_w[0] ;
 wire \clkgen.delay_155ns_1.genblk1[0].dly_binary.signal_w[1] ;
 wire \clkgen.delay_155ns_1.genblk1[1].dly_binary.bypass_in ;
 wire \clkgen.delay_155ns_1.genblk1[1].dly_binary.out ;
 wire \clkgen.delay_155ns_1.genblk1[1].dly_binary.signal_w[0] ;
 wire \clkgen.delay_155ns_1.genblk1[1].dly_binary.signal_w[1] ;
 wire \clkgen.delay_155ns_1.genblk1[1].dly_binary.signal_w[2] ;
 wire \clkgen.delay_155ns_1.genblk1[2].dly_binary.bypass_in ;
 wire \clkgen.delay_155ns_1.genblk1[2].dly_binary.out ;
 wire \clkgen.delay_155ns_1.genblk1[2].dly_binary.signal_w[0] ;
 wire \clkgen.delay_155ns_1.genblk1[2].dly_binary.signal_w[1] ;
 wire \clkgen.delay_155ns_1.genblk1[2].dly_binary.signal_w[2] ;
 wire \clkgen.delay_155ns_1.genblk1[2].dly_binary.signal_w[3] ;
 wire \clkgen.delay_155ns_1.genblk1[2].dly_binary.signal_w[4] ;
 wire \clkgen.delay_155ns_1.genblk1[3].dly_binary.bypass_in ;
 wire \clkgen.delay_155ns_1.genblk1[3].dly_binary.out ;
 wire \clkgen.delay_155ns_1.genblk1[3].dly_binary.signal_w[0] ;
 wire \clkgen.delay_155ns_1.genblk1[3].dly_binary.signal_w[1] ;
 wire \clkgen.delay_155ns_1.genblk1[3].dly_binary.signal_w[2] ;
 wire \clkgen.delay_155ns_1.genblk1[3].dly_binary.signal_w[3] ;
 wire \clkgen.delay_155ns_1.genblk1[3].dly_binary.signal_w[4] ;
 wire \clkgen.delay_155ns_1.genblk1[3].dly_binary.signal_w[5] ;
 wire \clkgen.delay_155ns_1.genblk1[3].dly_binary.signal_w[6] ;
 wire \clkgen.delay_155ns_1.genblk1[3].dly_binary.signal_w[7] ;
 wire \clkgen.delay_155ns_1.genblk1[3].dly_binary.signal_w[8] ;
 wire \clkgen.delay_155ns_1.genblk1[4].dly_binary.bypass_in ;
 wire \clkgen.delay_155ns_1.genblk1[4].dly_binary.out ;
 wire \clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[0] ;
 wire \clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[10] ;
 wire \clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[11] ;
 wire \clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[12] ;
 wire \clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[13] ;
 wire \clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[14] ;
 wire \clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[15] ;
 wire \clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[16] ;
 wire \clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[1] ;
 wire \clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[2] ;
 wire \clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[3] ;
 wire \clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[4] ;
 wire \clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[5] ;
 wire \clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[6] ;
 wire \clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[7] ;
 wire \clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[8] ;
 wire \clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[9] ;
 wire \clkgen.delay_155ns_2.bypass_enable_w[0] ;
 wire \clkgen.delay_155ns_2.bypass_enable_w[1] ;
 wire \clkgen.delay_155ns_2.bypass_enable_w[2] ;
 wire \clkgen.delay_155ns_2.bypass_enable_w[3] ;
 wire \clkgen.delay_155ns_2.bypass_enable_w[4] ;
 wire \clkgen.delay_155ns_2.enable_dlycontrol_w ;
 wire \clkgen.delay_155ns_2.genblk1[0].dly_binary.bypass_in ;
 wire \clkgen.delay_155ns_2.genblk1[0].dly_binary.out ;
 wire \clkgen.delay_155ns_2.genblk1[0].dly_binary.signal_w[0] ;
 wire \clkgen.delay_155ns_2.genblk1[0].dly_binary.signal_w[1] ;
 wire \clkgen.delay_155ns_2.genblk1[1].dly_binary.bypass_in ;
 wire \clkgen.delay_155ns_2.genblk1[1].dly_binary.out ;
 wire \clkgen.delay_155ns_2.genblk1[1].dly_binary.signal_w[0] ;
 wire \clkgen.delay_155ns_2.genblk1[1].dly_binary.signal_w[1] ;
 wire \clkgen.delay_155ns_2.genblk1[1].dly_binary.signal_w[2] ;
 wire \clkgen.delay_155ns_2.genblk1[2].dly_binary.bypass_in ;
 wire \clkgen.delay_155ns_2.genblk1[2].dly_binary.out ;
 wire \clkgen.delay_155ns_2.genblk1[2].dly_binary.signal_w[0] ;
 wire \clkgen.delay_155ns_2.genblk1[2].dly_binary.signal_w[1] ;
 wire \clkgen.delay_155ns_2.genblk1[2].dly_binary.signal_w[2] ;
 wire \clkgen.delay_155ns_2.genblk1[2].dly_binary.signal_w[3] ;
 wire \clkgen.delay_155ns_2.genblk1[2].dly_binary.signal_w[4] ;
 wire \clkgen.delay_155ns_2.genblk1[3].dly_binary.bypass_in ;
 wire \clkgen.delay_155ns_2.genblk1[3].dly_binary.out ;
 wire \clkgen.delay_155ns_2.genblk1[3].dly_binary.signal_w[0] ;
 wire \clkgen.delay_155ns_2.genblk1[3].dly_binary.signal_w[1] ;
 wire \clkgen.delay_155ns_2.genblk1[3].dly_binary.signal_w[2] ;
 wire \clkgen.delay_155ns_2.genblk1[3].dly_binary.signal_w[3] ;
 wire \clkgen.delay_155ns_2.genblk1[3].dly_binary.signal_w[4] ;
 wire \clkgen.delay_155ns_2.genblk1[3].dly_binary.signal_w[5] ;
 wire \clkgen.delay_155ns_2.genblk1[3].dly_binary.signal_w[6] ;
 wire \clkgen.delay_155ns_2.genblk1[3].dly_binary.signal_w[7] ;
 wire \clkgen.delay_155ns_2.genblk1[3].dly_binary.signal_w[8] ;
 wire \clkgen.delay_155ns_2.genblk1[4].dly_binary.bypass_in ;
 wire \clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[0] ;
 wire \clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[10] ;
 wire \clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[11] ;
 wire \clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[12] ;
 wire \clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[13] ;
 wire \clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[14] ;
 wire \clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[15] ;
 wire \clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[16] ;
 wire \clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[1] ;
 wire \clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[2] ;
 wire \clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[3] ;
 wire \clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[4] ;
 wire \clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[5] ;
 wire \clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[6] ;
 wire \clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[7] ;
 wire \clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[8] ;
 wire \clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[9] ;
 wire \clkgen.delay_155ns_3.bypass_enable_w[0] ;
 wire \clkgen.delay_155ns_3.bypass_enable_w[1] ;
 wire \clkgen.delay_155ns_3.bypass_enable_w[2] ;
 wire \clkgen.delay_155ns_3.bypass_enable_w[3] ;
 wire \clkgen.delay_155ns_3.bypass_enable_w[4] ;
 wire \clkgen.delay_155ns_3.enable_dlycontrol_w ;
 wire \clkgen.delay_155ns_3.genblk1[0].dly_binary.bypass_in ;
 wire \clkgen.delay_155ns_3.genblk1[0].dly_binary.in ;
 wire \clkgen.delay_155ns_3.genblk1[0].dly_binary.out ;
 wire \clkgen.delay_155ns_3.genblk1[0].dly_binary.signal_w[0] ;
 wire \clkgen.delay_155ns_3.genblk1[0].dly_binary.signal_w[1] ;
 wire \clkgen.delay_155ns_3.genblk1[1].dly_binary.bypass_in ;
 wire \clkgen.delay_155ns_3.genblk1[1].dly_binary.out ;
 wire \clkgen.delay_155ns_3.genblk1[1].dly_binary.signal_w[0] ;
 wire \clkgen.delay_155ns_3.genblk1[1].dly_binary.signal_w[1] ;
 wire \clkgen.delay_155ns_3.genblk1[1].dly_binary.signal_w[2] ;
 wire \clkgen.delay_155ns_3.genblk1[2].dly_binary.bypass_in ;
 wire \clkgen.delay_155ns_3.genblk1[2].dly_binary.out ;
 wire \clkgen.delay_155ns_3.genblk1[2].dly_binary.signal_w[0] ;
 wire \clkgen.delay_155ns_3.genblk1[2].dly_binary.signal_w[1] ;
 wire \clkgen.delay_155ns_3.genblk1[2].dly_binary.signal_w[2] ;
 wire \clkgen.delay_155ns_3.genblk1[2].dly_binary.signal_w[3] ;
 wire \clkgen.delay_155ns_3.genblk1[2].dly_binary.signal_w[4] ;
 wire \clkgen.delay_155ns_3.genblk1[3].dly_binary.bypass_in ;
 wire \clkgen.delay_155ns_3.genblk1[3].dly_binary.out ;
 wire \clkgen.delay_155ns_3.genblk1[3].dly_binary.signal_w[0] ;
 wire \clkgen.delay_155ns_3.genblk1[3].dly_binary.signal_w[1] ;
 wire \clkgen.delay_155ns_3.genblk1[3].dly_binary.signal_w[2] ;
 wire \clkgen.delay_155ns_3.genblk1[3].dly_binary.signal_w[3] ;
 wire \clkgen.delay_155ns_3.genblk1[3].dly_binary.signal_w[4] ;
 wire \clkgen.delay_155ns_3.genblk1[3].dly_binary.signal_w[5] ;
 wire \clkgen.delay_155ns_3.genblk1[3].dly_binary.signal_w[6] ;
 wire \clkgen.delay_155ns_3.genblk1[3].dly_binary.signal_w[7] ;
 wire \clkgen.delay_155ns_3.genblk1[3].dly_binary.signal_w[8] ;
 wire \clkgen.delay_155ns_3.genblk1[4].dly_binary.bypass_in ;
 wire \clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[0] ;
 wire \clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[10] ;
 wire \clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[11] ;
 wire \clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[12] ;
 wire \clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[13] ;
 wire \clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[14] ;
 wire \clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[15] ;
 wire \clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[16] ;
 wire \clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[1] ;
 wire \clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[2] ;
 wire \clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[3] ;
 wire \clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[4] ;
 wire \clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[5] ;
 wire \clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[6] ;
 wire \clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[7] ;
 wire \clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[8] ;
 wire \clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[9] ;
 wire \clkgen.enable_loop_in ;
 wire \edgedetect.dly_315ns_1.bypass_enable_w[0] ;
 wire \edgedetect.dly_315ns_1.bypass_enable_w[1] ;
 wire \edgedetect.dly_315ns_1.bypass_enable_w[2] ;
 wire \edgedetect.dly_315ns_1.bypass_enable_w[3] ;
 wire \edgedetect.dly_315ns_1.bypass_enable_w[4] ;
 wire \edgedetect.dly_315ns_1.bypass_enable_w[5] ;
 wire \edgedetect.dly_315ns_1.enable_dlycontrol_w ;
 wire \edgedetect.dly_315ns_1.genblk1[0].dly_binary.bypass_in ;
 wire \edgedetect.dly_315ns_1.genblk1[0].dly_binary.in ;
 wire \edgedetect.dly_315ns_1.genblk1[0].dly_binary.out ;
 wire \edgedetect.dly_315ns_1.genblk1[0].dly_binary.signal_w[0] ;
 wire \edgedetect.dly_315ns_1.genblk1[0].dly_binary.signal_w[1] ;
 wire \edgedetect.dly_315ns_1.genblk1[1].dly_binary.bypass_in ;
 wire \edgedetect.dly_315ns_1.genblk1[1].dly_binary.out ;
 wire \edgedetect.dly_315ns_1.genblk1[1].dly_binary.signal_w[0] ;
 wire \edgedetect.dly_315ns_1.genblk1[1].dly_binary.signal_w[1] ;
 wire \edgedetect.dly_315ns_1.genblk1[1].dly_binary.signal_w[2] ;
 wire \edgedetect.dly_315ns_1.genblk1[2].dly_binary.bypass_in ;
 wire \edgedetect.dly_315ns_1.genblk1[2].dly_binary.out ;
 wire \edgedetect.dly_315ns_1.genblk1[2].dly_binary.signal_w[0] ;
 wire \edgedetect.dly_315ns_1.genblk1[2].dly_binary.signal_w[1] ;
 wire \edgedetect.dly_315ns_1.genblk1[2].dly_binary.signal_w[2] ;
 wire \edgedetect.dly_315ns_1.genblk1[2].dly_binary.signal_w[3] ;
 wire \edgedetect.dly_315ns_1.genblk1[2].dly_binary.signal_w[4] ;
 wire \edgedetect.dly_315ns_1.genblk1[3].dly_binary.bypass_in ;
 wire \edgedetect.dly_315ns_1.genblk1[3].dly_binary.out ;
 wire \edgedetect.dly_315ns_1.genblk1[3].dly_binary.signal_w[0] ;
 wire \edgedetect.dly_315ns_1.genblk1[3].dly_binary.signal_w[1] ;
 wire \edgedetect.dly_315ns_1.genblk1[3].dly_binary.signal_w[2] ;
 wire \edgedetect.dly_315ns_1.genblk1[3].dly_binary.signal_w[3] ;
 wire \edgedetect.dly_315ns_1.genblk1[3].dly_binary.signal_w[4] ;
 wire \edgedetect.dly_315ns_1.genblk1[3].dly_binary.signal_w[5] ;
 wire \edgedetect.dly_315ns_1.genblk1[3].dly_binary.signal_w[6] ;
 wire \edgedetect.dly_315ns_1.genblk1[3].dly_binary.signal_w[7] ;
 wire \edgedetect.dly_315ns_1.genblk1[3].dly_binary.signal_w[8] ;
 wire \edgedetect.dly_315ns_1.genblk1[4].dly_binary.bypass_in ;
 wire \edgedetect.dly_315ns_1.genblk1[4].dly_binary.out ;
 wire \edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[0] ;
 wire \edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[10] ;
 wire \edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[11] ;
 wire \edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[12] ;
 wire \edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[13] ;
 wire \edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[14] ;
 wire \edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[15] ;
 wire \edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[16] ;
 wire \edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[1] ;
 wire \edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[2] ;
 wire \edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[3] ;
 wire \edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[4] ;
 wire \edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[5] ;
 wire \edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[6] ;
 wire \edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[7] ;
 wire \edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[8] ;
 wire \edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[9] ;
 wire \edgedetect.dly_315ns_1.genblk1[5].dly_binary.bypass_in ;
 wire \edgedetect.dly_315ns_1.genblk1[5].dly_binary.out ;
 wire \edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[0] ;
 wire \edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[10] ;
 wire \edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[11] ;
 wire \edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[12] ;
 wire \edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[13] ;
 wire \edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[14] ;
 wire \edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[15] ;
 wire \edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[16] ;
 wire \edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[17] ;
 wire \edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[18] ;
 wire \edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[19] ;
 wire \edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[1] ;
 wire \edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[20] ;
 wire \edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[21] ;
 wire \edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[22] ;
 wire \edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[23] ;
 wire \edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[24] ;
 wire \edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[25] ;
 wire \edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[26] ;
 wire \edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[27] ;
 wire \edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[28] ;
 wire \edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[29] ;
 wire \edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[2] ;
 wire \edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[30] ;
 wire \edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[31] ;
 wire \edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[32] ;
 wire \edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[3] ;
 wire \edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[4] ;
 wire \edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[5] ;
 wire \edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[6] ;
 wire \edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[7] ;
 wire \edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[8] ;
 wire \edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[9] ;
 wire \edgedetect.ena_in ;
 wire \edgedetect.start_conv_edge_w ;
 wire sample_n_1;
 wire sample_p_1;

 sky130_fd_sc_hd__diode_2 \ANTENNA_clkgen.delay_155ns_1.enablebuffer_A  (.DIODE(enable_dlycontrol_in),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkgen.delay_155ns_1.genblk1[0].control_invert_A  (.DIODE(dlycontrol1_in[0]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkgen.delay_155ns_1.genblk1[0].dly_binary.and_bypass_switch_A_N  (.DIODE(\clkgen.delay_155ns_1.genblk1[0].dly_binary.bypass_in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkgen.delay_155ns_1.genblk1[0].dly_binary.out_mux_S  (.DIODE(\clkgen.delay_155ns_1.genblk1[0].dly_binary.bypass_in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkgen.delay_155ns_1.genblk1[1].control_invert_A  (.DIODE(dlycontrol1_in[1]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkgen.delay_155ns_1.genblk1[2].control_invert_A  (.DIODE(dlycontrol1_in[2]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkgen.delay_155ns_1.genblk1[3].control_invert_A  (.DIODE(dlycontrol1_in[3]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkgen.delay_155ns_1.genblk1[3].dly_binary.and_bypass_switch_A_N  (.DIODE(\clkgen.delay_155ns_1.genblk1[3].dly_binary.bypass_in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkgen.delay_155ns_1.genblk1[3].dly_binary.out_mux_A0  (.DIODE(\clkgen.delay_155ns_1.genblk1[3].dly_binary.signal_w[8] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkgen.delay_155ns_1.genblk1[3].dly_binary.out_mux_S  (.DIODE(\clkgen.delay_155ns_1.genblk1[3].dly_binary.bypass_in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkgen.delay_155ns_1.genblk1[4].control_invert_A  (.DIODE(dlycontrol1_in[4]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkgen.delay_155ns_1.genblk1[4].dly_binary.and_bypass_switch_B  (.DIODE(\clkgen.delay_155ns_1.genblk1[3].dly_binary.out ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkgen.delay_155ns_1.genblk1[4].dly_binary.out_mux_A1  (.DIODE(\clkgen.delay_155ns_1.genblk1[3].dly_binary.out ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkgen.delay_155ns_2.enablebuffer_A  (.DIODE(enable_dlycontrol_in),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkgen.delay_155ns_2.genblk1[0].control_invert_A  (.DIODE(dlycontrol2_in[0]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkgen.delay_155ns_2.genblk1[0].dly_binary.and_bypass_switch_B  (.DIODE(\clkgen.clk_dig_out ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkgen.delay_155ns_2.genblk1[0].dly_binary.out_mux_A1  (.DIODE(\clkgen.clk_dig_out ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkgen.delay_155ns_2.genblk1[1].control_invert_A  (.DIODE(dlycontrol2_in[1]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkgen.delay_155ns_2.genblk1[1].dly_binary.and_bypass_switch_A_N  (.DIODE(\clkgen.delay_155ns_2.genblk1[1].dly_binary.bypass_in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkgen.delay_155ns_2.genblk1[1].dly_binary.and_bypass_switch_B  (.DIODE(\clkgen.delay_155ns_2.genblk1[0].dly_binary.out ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkgen.delay_155ns_2.genblk1[1].dly_binary.out_mux_A1  (.DIODE(\clkgen.delay_155ns_2.genblk1[0].dly_binary.out ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkgen.delay_155ns_2.genblk1[1].dly_binary.out_mux_S  (.DIODE(\clkgen.delay_155ns_2.genblk1[1].dly_binary.bypass_in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkgen.delay_155ns_2.genblk1[2].control_invert_A  (.DIODE(dlycontrol2_in[2]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkgen.delay_155ns_2.genblk1[2].dly_binary.and_bypass_switch_A_N  (.DIODE(\clkgen.delay_155ns_2.genblk1[2].dly_binary.bypass_in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkgen.delay_155ns_2.genblk1[2].dly_binary.out_mux_S  (.DIODE(\clkgen.delay_155ns_2.genblk1[2].dly_binary.bypass_in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkgen.delay_155ns_2.genblk1[3].control_invert_A  (.DIODE(dlycontrol2_in[3]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkgen.delay_155ns_2.genblk1[3].dly_binary.and_bypass_switch_A_N  (.DIODE(\clkgen.delay_155ns_2.genblk1[3].dly_binary.bypass_in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkgen.delay_155ns_2.genblk1[3].dly_binary.out_mux_S  (.DIODE(\clkgen.delay_155ns_2.genblk1[3].dly_binary.bypass_in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkgen.delay_155ns_2.genblk1[4].control_invert_A  (.DIODE(dlycontrol2_in[4]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkgen.delay_155ns_2.genblk1[4].dly_binary.and_bypass_switch_A_N  (.DIODE(\clkgen.delay_155ns_2.genblk1[4].dly_binary.bypass_in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkgen.delay_155ns_2.genblk1[4].dly_binary.out_mux_A0  (.DIODE(\clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[16] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkgen.delay_155ns_2.genblk1[4].dly_binary.out_mux_S  (.DIODE(\clkgen.delay_155ns_2.genblk1[4].dly_binary.bypass_in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkgen.delay_155ns_3.enablebuffer_A  (.DIODE(enable_dlycontrol_in),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkgen.delay_155ns_3.genblk1[0].control_invert_A  (.DIODE(dlycontrol3_in[0]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkgen.delay_155ns_3.genblk1[1].control_invert_A  (.DIODE(dlycontrol3_in[1]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkgen.delay_155ns_3.genblk1[2].control_invert_A  (.DIODE(dlycontrol3_in[2]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkgen.delay_155ns_3.genblk1[3].control_invert_A  (.DIODE(dlycontrol3_in[3]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkgen.delay_155ns_3.genblk1[4].control_invert_A  (.DIODE(dlycontrol3_in[4]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 ANTENNA_delay_sample_n12_in (.DIODE(sample_n_in),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 ANTENNA_delay_sample_p11_in (.DIODE(sample_p_in),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_edgedetect.dly_315ns_1.enablebuffer_A  (.DIODE(enable_dlycontrol_in),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_edgedetect.dly_315ns_1.genblk1[0].control_invert_A  (.DIODE(dlycontrol4_in[0]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_edgedetect.dly_315ns_1.genblk1[0].dly_binary.and_bypass_switch_A_N  (.DIODE(\edgedetect.dly_315ns_1.genblk1[0].dly_binary.bypass_in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_edgedetect.dly_315ns_1.genblk1[0].dly_binary.and_bypass_switch_B  (.DIODE(\edgedetect.dly_315ns_1.genblk1[0].dly_binary.in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_edgedetect.dly_315ns_1.genblk1[0].dly_binary.out_mux_A1  (.DIODE(\edgedetect.dly_315ns_1.genblk1[0].dly_binary.in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_edgedetect.dly_315ns_1.genblk1[0].dly_binary.out_mux_S  (.DIODE(\edgedetect.dly_315ns_1.genblk1[0].dly_binary.bypass_in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_edgedetect.dly_315ns_1.genblk1[1].control_invert_A  (.DIODE(dlycontrol4_in[1]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_edgedetect.dly_315ns_1.genblk1[1].dly_binary.and_bypass_switch_B  (.DIODE(\edgedetect.dly_315ns_1.genblk1[0].dly_binary.out ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_edgedetect.dly_315ns_1.genblk1[1].dly_binary.out_mux_A1  (.DIODE(\edgedetect.dly_315ns_1.genblk1[0].dly_binary.out ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_edgedetect.dly_315ns_1.genblk1[2].control_invert_A  (.DIODE(dlycontrol4_in[2]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_edgedetect.dly_315ns_1.genblk1[3].control_invert_A  (.DIODE(dlycontrol4_in[3]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_edgedetect.dly_315ns_1.genblk1[3].dly_binary.genblk1[0].delay_unit_in  (.DIODE(\edgedetect.dly_315ns_1.genblk1[3].dly_binary.signal_w[0] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_edgedetect.dly_315ns_1.genblk1[4].control_invert_A  (.DIODE(dlycontrol4_in[4]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_edgedetect.dly_315ns_1.genblk1[4].dly_binary.genblk1[0].delay_unit_in  (.DIODE(\edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[0] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_edgedetect.dly_315ns_1.genblk1[5].control_invert_A  (.DIODE(dlycontrol4_in[5]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_edgedetect.nor1_B_N  (.DIODE(\edgedetect.dly_315ns_1.genblk1[0].dly_binary.in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_edgedetect.or1_A  (.DIODE(\edgedetect.start_conv_edge_w ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 \ANTENNA_edgedetect.or1_B  (.DIODE(\edgedetect.ena_in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 ANTENNA_inbuf_1_A (.DIODE(ena_in),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 ANTENNA_inbuf_2_A (.DIODE(start_conv_in),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 ANTENNA_inbuf_3_A (.DIODE(ndecision_finish_in),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__diode_2 ANTENNA_outbuf_1_A (.DIODE(\clkgen.clk_dig_out ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_0_122 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_0_125 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_0_136 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_0_146 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_0_153 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_0_156 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_0_182 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_0_187 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_0_194 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_0_203 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_0_210 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_0_216 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_0_218 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_0_223 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_0_229 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_0_235 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_0_241 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_0_247 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_0_249 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_0_253 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_0_259 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_265 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_0_277 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_280 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_0_29 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_292 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_0_3 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_0_304 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_311 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_0_32 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_0_323 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_0_335 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_0_342 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_0_60 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_0_63 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_0_91 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_0_94 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_100 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_10_125 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_10_153 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_10_156 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_10_16 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_10_164 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_10_174 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_182 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_10_207 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_10_214 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_10_218 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_10_244 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_252 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_10_277 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_10_280 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_10_284 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_10_29 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_292 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_10_3 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_10_317 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_10_32 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_10_323 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_10_335 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_10_342 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_10_58 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_10_66 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_10_91 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_10_94 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_11_122 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_11_125 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_11_151 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_11_179 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_185 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_11_187 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_11_19 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_11_213 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_11_241 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_247 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_11_249 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_11_256 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_11_263 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_11_270 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_11_276 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_11_282 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_11_288 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_11_294 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_11_3 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_11_300 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_11_306 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_11_311 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_315 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_11_32 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_11_327 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_11_339 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_343 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_11_60 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_11_63 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_11_89 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_9 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_11_97 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_12_10 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_12_104 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_12_117 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_12_145 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_12_152 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_12_156 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_12_164 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_172 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_12_197 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_12_207 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_12_214 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_12_218 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_12_226 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_232 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_12_257 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_12_266 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_12_273 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_12_280 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_12_284 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_12_29 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_12_290 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_12_296 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_12_3 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_12_302 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_12_308 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_12_314 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_12_32 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_12_320 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_12_326 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_12_338 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_12_342 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_12_38 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_12_63 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_12_91 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_12_94 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_13_113 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_13_122 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_13_125 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_13_133 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_13_161 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_13_174 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_13_184 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_13_187 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_13_195 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_13_227 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_13_236 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_13_245 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_13_249 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_13_275 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_13_282 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_13_288 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_13_294 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_13_3 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_13_300 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_13_306 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_13_31 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_13_311 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_317 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_13_342 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_13_59 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_13_63 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_13_74 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_13_84 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_13_88 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_100 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_14_125 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_14_153 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_14_156 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_160 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_14_185 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_14_213 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_14_218 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_14_244 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_14_272 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_278 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_14_280 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_14_29 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_14_3 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_14_306 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_314 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_14_32 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_14_339 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_14_342 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_14_38 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_14_63 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_14_91 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_14_94 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_15_116 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_15_122 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_15_125 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_131 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_15_156 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_15_184 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_15_187 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_191 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_15_216 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_15_246 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_15_249 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_15_256 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_15_284 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_15_29 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_15_291 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_15_298 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_15_3 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_15_304 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_15_311 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_15_337 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_343 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_15_59 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_15_63 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_15_74 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_15_87 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_15_91 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_100 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_16_125 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_16_153 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_16_156 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_16_167 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_173 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_16_198 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_16_208 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_16_215 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_16_218 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_16_244 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_252 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_16_277 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_16_280 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_16_29 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_16_3 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_16_306 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_16_32 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_16_334 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_340 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_16_342 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_16_38 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_16_63 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_16_91 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_16_94 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_17_122 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_17_125 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_131 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_156 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_17_184 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_17_187 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_198 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_202 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_227 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_237 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_17_246 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_17_249 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_275 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_3 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_17_303 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_309 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_17_311 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_32 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_17_337 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_343 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_17_60 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_17_63 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_69 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_17_7 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_17_94 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_18_100 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_125 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_18_153 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_156 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_18_160 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_185 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_213 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_18_218 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_244 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_18_272 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_18_278 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_18_280 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_284 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_18_29 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_18_3 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_312 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_318 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_18_32 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_18_324 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_336 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_18_340 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_18_342 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_18_38 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_18_63 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_18_91 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_18_94 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_120 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_19_125 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_151 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_19_156 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_182 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_19_187 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_213 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_19_218 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_244 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_19_249 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_256 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_265 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_274 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_19_278 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_19_280 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_285 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_19_29 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_292 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_298 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_19_3 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_19_304 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_19_311 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_315 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_32 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_19_327 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_19_339 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_19_342 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_19_60 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_19_63 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_19_91 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_19_94 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_1_122 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_1_125 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_1_153 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_159 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_1_184 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_1_187 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_193 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_1_218 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_1_225 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_1_231 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_1_237 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_1_243 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_247 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_1_249 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_1_253 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_259 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_271 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_283 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_295 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_1_3 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_1_307 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_311 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_1_32 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_1_323 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_1_335 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_343 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_1_60 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_1_63 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_69 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_1_7 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_1_94 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_100 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_2_125 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_2_153 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_2_156 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_2_164 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_2_174 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_2_206 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_2_215 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_2_218 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_2_223 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_2_230 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_2_237 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_2_243 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_2_249 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_2_255 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_2_261 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_2_267 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_2_273 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_280 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_2_29 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_292 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_2_3 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_304 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_316 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_2_32 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_2_328 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_340 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_2_342 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_2_38 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_2_63 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_2_91 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_2_94 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_3_122 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_3_125 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_3_151 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_3_181 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_185 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_3_187 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_3_213 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_3_223 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_3_232 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_3_239 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_3_246 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_3_249 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_3_253 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_3_259 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_3_265 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_3_271 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_3_277 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_283 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_295 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_3_3 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_3_30 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_3_307 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_311 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_3_323 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_3_335 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_343 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_3_60 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_3_63 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_3_69 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_3_94 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_100 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_4_125 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_4_153 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_4_156 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_4_167 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_4_173 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_4_201 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_4_211 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_4_218 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_4_226 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_4_235 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_4_242 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_4_249 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_4_256 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_4_262 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_4_268 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_4_274 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_278 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_4_280 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_4_284 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_4_29 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_290 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_4_3 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_302 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_314 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_4_32 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_4_326 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_4_338 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_4_342 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_4_38 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_4_63 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_4_91 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_4_94 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_5_110 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_114 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_5_121 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_5_125 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_5_13 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_5_142 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_5_174 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_5_184 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_5_187 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_5_213 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_5_222 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_5_231 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_5_240 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_5_246 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_5_249 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_253 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_5_278 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_5_284 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_290 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_5_3 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_5_302 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_311 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_5_32 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_ef_sc_hd__decap_12 FILLER_5_323 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_5_335 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_343 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_5_60 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_5_63 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_5_68 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_5_81 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_5_85 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_6_120 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_128 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_6_153 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_6_156 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_162 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_6_187 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_6_215 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_6_218 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_6_244 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_6_272 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_278 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_6_280 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_6_29 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_6_3 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_6_306 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_6_32 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_6_334 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_340 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_6_342 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_6_43 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_6_47 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_6_57 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_6_85 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_6_91 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_6_94 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_7_122 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_7_125 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_131 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_7_156 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_7_184 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_7_187 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_7_195 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_203 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_7_228 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_7_237 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_7_246 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_7_249 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_7_275 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_7_3 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_7_303 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_309 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_7_311 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_7_32 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_7_337 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_343 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_7_60 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_7_63 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_69 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_7_7 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_7_94 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_8_10 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_8_120 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_128 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_8_153 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_8_156 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_8_167 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_8_177 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_181 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_8_206 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_8_215 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_8_218 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_8_244 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_8_272 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_278 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_8_280 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_8_29 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_8_3 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_8_306 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_314 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 FILLER_8_32 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_8_339 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_8_342 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_8_44 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_50 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_8_75 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_8_88 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_8_92 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_8_94 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_9_122 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_9_125 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_8 FILLER_9_151 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_159 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_9_184 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_9_187 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_9_19 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_9_195 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_9_223 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_9_233 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_9_242 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_9_249 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_9_275 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_9_3 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_9_303 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_309 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_9_311 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_9_32 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_9_337 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_343 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_2 FILLER_9_60 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_4 FILLER_9_63 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_9 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_6 FILLER_9_91 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__fill_1 FILLER_9_97 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_0 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_1 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_10 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_11 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_12 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_13 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_14 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_15 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_16 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_17 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_18 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_19 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_2 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_20 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_21 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_22 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_23 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_24 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_25 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_26 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_27 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_28 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_29 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_3 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_30 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_31 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_32 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_33 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_34 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_35 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_36 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_37 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_38 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_39 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_4 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_5 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_6 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_7 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_8 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__decap_3 PHY_9 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_40 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_41 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_42 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_43 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_44 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_45 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_46 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_47 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_48 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_49 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_50 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_51 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_52 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_53 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_54 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_55 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_56 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_57 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_58 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_59 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_60 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_61 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_62 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_63 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_64 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_65 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_66 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_67 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_68 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_69 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_70 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_71 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_72 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_73 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_74 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_75 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_76 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_77 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_78 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_79 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_80 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_81 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_82 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_83 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_84 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_85 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_86 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_87 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_88 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_89 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_90 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_91 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_92 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_93 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_94 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_95 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_96 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_97 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 (.VGND(VSS),
    .VPWR(VDD));
 sky130_fd_sc_hd__inv_2 \clkgen.clkdig_inverter  (.A(\clkgen.delay_155ns_1.genblk1[4].dly_binary.out ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(\clkgen.clk_dig_out ));
 sky130_fd_sc_hd__buf_4 \clkgen.delay_155ns_1.enablebuffer  (.A(enable_dlycontrol_in),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_1.enable_dlycontrol_w ));
 sky130_fd_sc_hd__and2_1 \clkgen.delay_155ns_1.genblk1[0].bypass_enable  (.A(\clkgen.delay_155ns_1.enable_dlycontrol_w ),
    .B(\clkgen.delay_155ns_1.bypass_enable_w[0] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_1.genblk1[0].dly_binary.bypass_in ));
 sky130_fd_sc_hd__inv_2 \clkgen.delay_155ns_1.genblk1[0].control_invert  (.A(dlycontrol1_in[0]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(\clkgen.delay_155ns_1.bypass_enable_w[0] ));
 sky130_fd_sc_hd__and2b_1 \clkgen.delay_155ns_1.genblk1[0].dly_binary.and_bypass_switch  (.A_N(\clkgen.delay_155ns_1.genblk1[0].dly_binary.bypass_in ),
    .B(\clkgen.delay_155ns_1.genblk1[0].dly_binary.in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_1.genblk1[0].dly_binary.signal_w[0] ));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_1.genblk1[0].dly_binary.genblk1[0].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_1.genblk1[0].dly_binary.signal_w[0] ),
    .out(\clkgen.delay_155ns_1.genblk1[0].dly_binary.signal_w[1] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_fd_sc_hd__mux2_1 \clkgen.delay_155ns_1.genblk1[0].dly_binary.out_mux  (.A0(\clkgen.delay_155ns_1.genblk1[0].dly_binary.signal_w[1] ),
    .A1(\clkgen.delay_155ns_1.genblk1[0].dly_binary.in ),
    .S(\clkgen.delay_155ns_1.genblk1[0].dly_binary.bypass_in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_1.genblk1[0].dly_binary.out ));
 sky130_fd_sc_hd__and2_1 \clkgen.delay_155ns_1.genblk1[1].bypass_enable  (.A(\clkgen.delay_155ns_1.enable_dlycontrol_w ),
    .B(\clkgen.delay_155ns_1.bypass_enable_w[1] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_1.genblk1[1].dly_binary.bypass_in ));
 sky130_fd_sc_hd__inv_2 \clkgen.delay_155ns_1.genblk1[1].control_invert  (.A(dlycontrol1_in[1]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(\clkgen.delay_155ns_1.bypass_enable_w[1] ));
 sky130_fd_sc_hd__and2b_1 \clkgen.delay_155ns_1.genblk1[1].dly_binary.and_bypass_switch  (.A_N(\clkgen.delay_155ns_1.genblk1[1].dly_binary.bypass_in ),
    .B(\clkgen.delay_155ns_1.genblk1[0].dly_binary.out ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_1.genblk1[1].dly_binary.signal_w[0] ));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_1.genblk1[1].dly_binary.genblk1[0].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_1.genblk1[1].dly_binary.signal_w[0] ),
    .out(\clkgen.delay_155ns_1.genblk1[1].dly_binary.signal_w[1] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_1.genblk1[1].dly_binary.genblk1[1].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_1.genblk1[1].dly_binary.signal_w[1] ),
    .out(\clkgen.delay_155ns_1.genblk1[1].dly_binary.signal_w[2] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_fd_sc_hd__mux2_1 \clkgen.delay_155ns_1.genblk1[1].dly_binary.out_mux  (.A0(\clkgen.delay_155ns_1.genblk1[1].dly_binary.signal_w[2] ),
    .A1(\clkgen.delay_155ns_1.genblk1[0].dly_binary.out ),
    .S(\clkgen.delay_155ns_1.genblk1[1].dly_binary.bypass_in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_1.genblk1[1].dly_binary.out ));
 sky130_fd_sc_hd__and2_1 \clkgen.delay_155ns_1.genblk1[2].bypass_enable  (.A(\clkgen.delay_155ns_1.enable_dlycontrol_w ),
    .B(\clkgen.delay_155ns_1.bypass_enable_w[2] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_1.genblk1[2].dly_binary.bypass_in ));
 sky130_fd_sc_hd__inv_2 \clkgen.delay_155ns_1.genblk1[2].control_invert  (.A(dlycontrol1_in[2]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(\clkgen.delay_155ns_1.bypass_enable_w[2] ));
 sky130_fd_sc_hd__and2b_1 \clkgen.delay_155ns_1.genblk1[2].dly_binary.and_bypass_switch  (.A_N(\clkgen.delay_155ns_1.genblk1[2].dly_binary.bypass_in ),
    .B(\clkgen.delay_155ns_1.genblk1[1].dly_binary.out ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_1.genblk1[2].dly_binary.signal_w[0] ));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_1.genblk1[2].dly_binary.genblk1[0].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_1.genblk1[2].dly_binary.signal_w[0] ),
    .out(\clkgen.delay_155ns_1.genblk1[2].dly_binary.signal_w[1] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_1.genblk1[2].dly_binary.genblk1[1].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_1.genblk1[2].dly_binary.signal_w[1] ),
    .out(\clkgen.delay_155ns_1.genblk1[2].dly_binary.signal_w[2] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_1.genblk1[2].dly_binary.genblk1[2].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_1.genblk1[2].dly_binary.signal_w[2] ),
    .out(\clkgen.delay_155ns_1.genblk1[2].dly_binary.signal_w[3] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_1.genblk1[2].dly_binary.genblk1[3].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_1.genblk1[2].dly_binary.signal_w[3] ),
    .out(\clkgen.delay_155ns_1.genblk1[2].dly_binary.signal_w[4] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_fd_sc_hd__mux2_1 \clkgen.delay_155ns_1.genblk1[2].dly_binary.out_mux  (.A0(\clkgen.delay_155ns_1.genblk1[2].dly_binary.signal_w[4] ),
    .A1(\clkgen.delay_155ns_1.genblk1[1].dly_binary.out ),
    .S(\clkgen.delay_155ns_1.genblk1[2].dly_binary.bypass_in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_1.genblk1[2].dly_binary.out ));
 sky130_fd_sc_hd__and2_1 \clkgen.delay_155ns_1.genblk1[3].bypass_enable  (.A(\clkgen.delay_155ns_1.enable_dlycontrol_w ),
    .B(\clkgen.delay_155ns_1.bypass_enable_w[3] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_1.genblk1[3].dly_binary.bypass_in ));
 sky130_fd_sc_hd__inv_2 \clkgen.delay_155ns_1.genblk1[3].control_invert  (.A(dlycontrol1_in[3]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(\clkgen.delay_155ns_1.bypass_enable_w[3] ));
 sky130_fd_sc_hd__and2b_1 \clkgen.delay_155ns_1.genblk1[3].dly_binary.and_bypass_switch  (.A_N(\clkgen.delay_155ns_1.genblk1[3].dly_binary.bypass_in ),
    .B(\clkgen.delay_155ns_1.genblk1[2].dly_binary.out ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_1.genblk1[3].dly_binary.signal_w[0] ));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_1.genblk1[3].dly_binary.genblk1[0].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_1.genblk1[3].dly_binary.signal_w[0] ),
    .out(\clkgen.delay_155ns_1.genblk1[3].dly_binary.signal_w[1] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_1.genblk1[3].dly_binary.genblk1[1].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_1.genblk1[3].dly_binary.signal_w[1] ),
    .out(\clkgen.delay_155ns_1.genblk1[3].dly_binary.signal_w[2] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_1.genblk1[3].dly_binary.genblk1[2].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_1.genblk1[3].dly_binary.signal_w[2] ),
    .out(\clkgen.delay_155ns_1.genblk1[3].dly_binary.signal_w[3] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_1.genblk1[3].dly_binary.genblk1[3].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_1.genblk1[3].dly_binary.signal_w[3] ),
    .out(\clkgen.delay_155ns_1.genblk1[3].dly_binary.signal_w[4] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_1.genblk1[3].dly_binary.genblk1[4].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_1.genblk1[3].dly_binary.signal_w[4] ),
    .out(\clkgen.delay_155ns_1.genblk1[3].dly_binary.signal_w[5] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_1.genblk1[3].dly_binary.genblk1[5].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_1.genblk1[3].dly_binary.signal_w[5] ),
    .out(\clkgen.delay_155ns_1.genblk1[3].dly_binary.signal_w[6] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_1.genblk1[3].dly_binary.genblk1[6].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_1.genblk1[3].dly_binary.signal_w[6] ),
    .out(\clkgen.delay_155ns_1.genblk1[3].dly_binary.signal_w[7] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_1.genblk1[3].dly_binary.genblk1[7].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_1.genblk1[3].dly_binary.signal_w[7] ),
    .out(\clkgen.delay_155ns_1.genblk1[3].dly_binary.signal_w[8] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_fd_sc_hd__mux2_1 \clkgen.delay_155ns_1.genblk1[3].dly_binary.out_mux  (.A0(\clkgen.delay_155ns_1.genblk1[3].dly_binary.signal_w[8] ),
    .A1(\clkgen.delay_155ns_1.genblk1[2].dly_binary.out ),
    .S(\clkgen.delay_155ns_1.genblk1[3].dly_binary.bypass_in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_1.genblk1[3].dly_binary.out ));
 sky130_fd_sc_hd__and2_1 \clkgen.delay_155ns_1.genblk1[4].bypass_enable  (.A(\clkgen.delay_155ns_1.enable_dlycontrol_w ),
    .B(\clkgen.delay_155ns_1.bypass_enable_w[4] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_1.genblk1[4].dly_binary.bypass_in ));
 sky130_fd_sc_hd__inv_2 \clkgen.delay_155ns_1.genblk1[4].control_invert  (.A(dlycontrol1_in[4]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(\clkgen.delay_155ns_1.bypass_enable_w[4] ));
 sky130_fd_sc_hd__and2b_1 \clkgen.delay_155ns_1.genblk1[4].dly_binary.and_bypass_switch  (.A_N(\clkgen.delay_155ns_1.genblk1[4].dly_binary.bypass_in ),
    .B(\clkgen.delay_155ns_1.genblk1[3].dly_binary.out ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[0] ));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_1.genblk1[4].dly_binary.genblk1[0].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[0] ),
    .out(\clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[1] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_1.genblk1[4].dly_binary.genblk1[10].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[10] ),
    .out(\clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[11] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_1.genblk1[4].dly_binary.genblk1[11].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[11] ),
    .out(\clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[12] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_1.genblk1[4].dly_binary.genblk1[12].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[12] ),
    .out(\clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[13] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_1.genblk1[4].dly_binary.genblk1[13].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[13] ),
    .out(\clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[14] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_1.genblk1[4].dly_binary.genblk1[14].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[14] ),
    .out(\clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[15] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_1.genblk1[4].dly_binary.genblk1[15].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[15] ),
    .out(\clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[16] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_1.genblk1[4].dly_binary.genblk1[1].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[1] ),
    .out(\clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[2] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_1.genblk1[4].dly_binary.genblk1[2].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[2] ),
    .out(\clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[3] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_1.genblk1[4].dly_binary.genblk1[3].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[3] ),
    .out(\clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[4] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_1.genblk1[4].dly_binary.genblk1[4].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[4] ),
    .out(\clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[5] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_1.genblk1[4].dly_binary.genblk1[5].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[5] ),
    .out(\clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[6] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_1.genblk1[4].dly_binary.genblk1[6].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[6] ),
    .out(\clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[7] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_1.genblk1[4].dly_binary.genblk1[7].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[7] ),
    .out(\clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[8] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_1.genblk1[4].dly_binary.genblk1[8].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[8] ),
    .out(\clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[9] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_1.genblk1[4].dly_binary.genblk1[9].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[9] ),
    .out(\clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[10] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_fd_sc_hd__mux2_1 \clkgen.delay_155ns_1.genblk1[4].dly_binary.out_mux  (.A0(\clkgen.delay_155ns_1.genblk1[4].dly_binary.signal_w[16] ),
    .A1(\clkgen.delay_155ns_1.genblk1[3].dly_binary.out ),
    .S(\clkgen.delay_155ns_1.genblk1[4].dly_binary.bypass_in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_1.genblk1[4].dly_binary.out ));
 sky130_fd_sc_hd__buf_4 \clkgen.delay_155ns_2.enablebuffer  (.A(enable_dlycontrol_in),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_2.enable_dlycontrol_w ));
 sky130_fd_sc_hd__and2_1 \clkgen.delay_155ns_2.genblk1[0].bypass_enable  (.A(\clkgen.delay_155ns_2.enable_dlycontrol_w ),
    .B(\clkgen.delay_155ns_2.bypass_enable_w[0] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_2.genblk1[0].dly_binary.bypass_in ));
 sky130_fd_sc_hd__inv_2 \clkgen.delay_155ns_2.genblk1[0].control_invert  (.A(dlycontrol2_in[0]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(\clkgen.delay_155ns_2.bypass_enable_w[0] ));
 sky130_fd_sc_hd__and2b_1 \clkgen.delay_155ns_2.genblk1[0].dly_binary.and_bypass_switch  (.A_N(\clkgen.delay_155ns_2.genblk1[0].dly_binary.bypass_in ),
    .B(\clkgen.clk_dig_out ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_2.genblk1[0].dly_binary.signal_w[0] ));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_2.genblk1[0].dly_binary.genblk1[0].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_2.genblk1[0].dly_binary.signal_w[0] ),
    .out(\clkgen.delay_155ns_2.genblk1[0].dly_binary.signal_w[1] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_fd_sc_hd__mux2_1 \clkgen.delay_155ns_2.genblk1[0].dly_binary.out_mux  (.A0(\clkgen.delay_155ns_2.genblk1[0].dly_binary.signal_w[1] ),
    .A1(\clkgen.clk_dig_out ),
    .S(\clkgen.delay_155ns_2.genblk1[0].dly_binary.bypass_in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_2.genblk1[0].dly_binary.out ));
 sky130_fd_sc_hd__and2_1 \clkgen.delay_155ns_2.genblk1[1].bypass_enable  (.A(\clkgen.delay_155ns_2.enable_dlycontrol_w ),
    .B(\clkgen.delay_155ns_2.bypass_enable_w[1] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_2.genblk1[1].dly_binary.bypass_in ));
 sky130_fd_sc_hd__inv_2 \clkgen.delay_155ns_2.genblk1[1].control_invert  (.A(dlycontrol2_in[1]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(\clkgen.delay_155ns_2.bypass_enable_w[1] ));
 sky130_fd_sc_hd__and2b_1 \clkgen.delay_155ns_2.genblk1[1].dly_binary.and_bypass_switch  (.A_N(\clkgen.delay_155ns_2.genblk1[1].dly_binary.bypass_in ),
    .B(\clkgen.delay_155ns_2.genblk1[0].dly_binary.out ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_2.genblk1[1].dly_binary.signal_w[0] ));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_2.genblk1[1].dly_binary.genblk1[0].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_2.genblk1[1].dly_binary.signal_w[0] ),
    .out(\clkgen.delay_155ns_2.genblk1[1].dly_binary.signal_w[1] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_2.genblk1[1].dly_binary.genblk1[1].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_2.genblk1[1].dly_binary.signal_w[1] ),
    .out(\clkgen.delay_155ns_2.genblk1[1].dly_binary.signal_w[2] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_fd_sc_hd__mux2_1 \clkgen.delay_155ns_2.genblk1[1].dly_binary.out_mux  (.A0(\clkgen.delay_155ns_2.genblk1[1].dly_binary.signal_w[2] ),
    .A1(\clkgen.delay_155ns_2.genblk1[0].dly_binary.out ),
    .S(\clkgen.delay_155ns_2.genblk1[1].dly_binary.bypass_in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_2.genblk1[1].dly_binary.out ));
 sky130_fd_sc_hd__and2_1 \clkgen.delay_155ns_2.genblk1[2].bypass_enable  (.A(\clkgen.delay_155ns_2.enable_dlycontrol_w ),
    .B(\clkgen.delay_155ns_2.bypass_enable_w[2] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_2.genblk1[2].dly_binary.bypass_in ));
 sky130_fd_sc_hd__inv_2 \clkgen.delay_155ns_2.genblk1[2].control_invert  (.A(dlycontrol2_in[2]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(\clkgen.delay_155ns_2.bypass_enable_w[2] ));
 sky130_fd_sc_hd__and2b_1 \clkgen.delay_155ns_2.genblk1[2].dly_binary.and_bypass_switch  (.A_N(\clkgen.delay_155ns_2.genblk1[2].dly_binary.bypass_in ),
    .B(\clkgen.delay_155ns_2.genblk1[1].dly_binary.out ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_2.genblk1[2].dly_binary.signal_w[0] ));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_2.genblk1[2].dly_binary.genblk1[0].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_2.genblk1[2].dly_binary.signal_w[0] ),
    .out(\clkgen.delay_155ns_2.genblk1[2].dly_binary.signal_w[1] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_2.genblk1[2].dly_binary.genblk1[1].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_2.genblk1[2].dly_binary.signal_w[1] ),
    .out(\clkgen.delay_155ns_2.genblk1[2].dly_binary.signal_w[2] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_2.genblk1[2].dly_binary.genblk1[2].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_2.genblk1[2].dly_binary.signal_w[2] ),
    .out(\clkgen.delay_155ns_2.genblk1[2].dly_binary.signal_w[3] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_2.genblk1[2].dly_binary.genblk1[3].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_2.genblk1[2].dly_binary.signal_w[3] ),
    .out(\clkgen.delay_155ns_2.genblk1[2].dly_binary.signal_w[4] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_fd_sc_hd__mux2_1 \clkgen.delay_155ns_2.genblk1[2].dly_binary.out_mux  (.A0(\clkgen.delay_155ns_2.genblk1[2].dly_binary.signal_w[4] ),
    .A1(\clkgen.delay_155ns_2.genblk1[1].dly_binary.out ),
    .S(\clkgen.delay_155ns_2.genblk1[2].dly_binary.bypass_in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_2.genblk1[2].dly_binary.out ));
 sky130_fd_sc_hd__and2_1 \clkgen.delay_155ns_2.genblk1[3].bypass_enable  (.A(\clkgen.delay_155ns_2.enable_dlycontrol_w ),
    .B(\clkgen.delay_155ns_2.bypass_enable_w[3] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_2.genblk1[3].dly_binary.bypass_in ));
 sky130_fd_sc_hd__inv_2 \clkgen.delay_155ns_2.genblk1[3].control_invert  (.A(dlycontrol2_in[3]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(\clkgen.delay_155ns_2.bypass_enable_w[3] ));
 sky130_fd_sc_hd__and2b_1 \clkgen.delay_155ns_2.genblk1[3].dly_binary.and_bypass_switch  (.A_N(\clkgen.delay_155ns_2.genblk1[3].dly_binary.bypass_in ),
    .B(\clkgen.delay_155ns_2.genblk1[2].dly_binary.out ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_2.genblk1[3].dly_binary.signal_w[0] ));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_2.genblk1[3].dly_binary.genblk1[0].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_2.genblk1[3].dly_binary.signal_w[0] ),
    .out(\clkgen.delay_155ns_2.genblk1[3].dly_binary.signal_w[1] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_2.genblk1[3].dly_binary.genblk1[1].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_2.genblk1[3].dly_binary.signal_w[1] ),
    .out(\clkgen.delay_155ns_2.genblk1[3].dly_binary.signal_w[2] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_2.genblk1[3].dly_binary.genblk1[2].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_2.genblk1[3].dly_binary.signal_w[2] ),
    .out(\clkgen.delay_155ns_2.genblk1[3].dly_binary.signal_w[3] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_2.genblk1[3].dly_binary.genblk1[3].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_2.genblk1[3].dly_binary.signal_w[3] ),
    .out(\clkgen.delay_155ns_2.genblk1[3].dly_binary.signal_w[4] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_2.genblk1[3].dly_binary.genblk1[4].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_2.genblk1[3].dly_binary.signal_w[4] ),
    .out(\clkgen.delay_155ns_2.genblk1[3].dly_binary.signal_w[5] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_2.genblk1[3].dly_binary.genblk1[5].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_2.genblk1[3].dly_binary.signal_w[5] ),
    .out(\clkgen.delay_155ns_2.genblk1[3].dly_binary.signal_w[6] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_2.genblk1[3].dly_binary.genblk1[6].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_2.genblk1[3].dly_binary.signal_w[6] ),
    .out(\clkgen.delay_155ns_2.genblk1[3].dly_binary.signal_w[7] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_2.genblk1[3].dly_binary.genblk1[7].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_2.genblk1[3].dly_binary.signal_w[7] ),
    .out(\clkgen.delay_155ns_2.genblk1[3].dly_binary.signal_w[8] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_fd_sc_hd__mux2_1 \clkgen.delay_155ns_2.genblk1[3].dly_binary.out_mux  (.A0(\clkgen.delay_155ns_2.genblk1[3].dly_binary.signal_w[8] ),
    .A1(\clkgen.delay_155ns_2.genblk1[2].dly_binary.out ),
    .S(\clkgen.delay_155ns_2.genblk1[3].dly_binary.bypass_in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_2.genblk1[3].dly_binary.out ));
 sky130_fd_sc_hd__and2_1 \clkgen.delay_155ns_2.genblk1[4].bypass_enable  (.A(\clkgen.delay_155ns_2.enable_dlycontrol_w ),
    .B(\clkgen.delay_155ns_2.bypass_enable_w[4] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_2.genblk1[4].dly_binary.bypass_in ));
 sky130_fd_sc_hd__inv_2 \clkgen.delay_155ns_2.genblk1[4].control_invert  (.A(dlycontrol2_in[4]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(\clkgen.delay_155ns_2.bypass_enable_w[4] ));
 sky130_fd_sc_hd__and2b_1 \clkgen.delay_155ns_2.genblk1[4].dly_binary.and_bypass_switch  (.A_N(\clkgen.delay_155ns_2.genblk1[4].dly_binary.bypass_in ),
    .B(\clkgen.delay_155ns_2.genblk1[3].dly_binary.out ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[0] ));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_2.genblk1[4].dly_binary.genblk1[0].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[0] ),
    .out(\clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[1] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_2.genblk1[4].dly_binary.genblk1[10].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[10] ),
    .out(\clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[11] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_2.genblk1[4].dly_binary.genblk1[11].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[11] ),
    .out(\clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[12] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_2.genblk1[4].dly_binary.genblk1[12].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[12] ),
    .out(\clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[13] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_2.genblk1[4].dly_binary.genblk1[13].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[13] ),
    .out(\clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[14] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_2.genblk1[4].dly_binary.genblk1[14].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[14] ),
    .out(\clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[15] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_2.genblk1[4].dly_binary.genblk1[15].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[15] ),
    .out(\clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[16] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_2.genblk1[4].dly_binary.genblk1[1].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[1] ),
    .out(\clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[2] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_2.genblk1[4].dly_binary.genblk1[2].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[2] ),
    .out(\clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[3] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_2.genblk1[4].dly_binary.genblk1[3].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[3] ),
    .out(\clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[4] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_2.genblk1[4].dly_binary.genblk1[4].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[4] ),
    .out(\clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[5] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_2.genblk1[4].dly_binary.genblk1[5].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[5] ),
    .out(\clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[6] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_2.genblk1[4].dly_binary.genblk1[6].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[6] ),
    .out(\clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[7] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_2.genblk1[4].dly_binary.genblk1[7].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[7] ),
    .out(\clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[8] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_2.genblk1[4].dly_binary.genblk1[8].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[8] ),
    .out(\clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[9] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_2.genblk1[4].dly_binary.genblk1[9].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[9] ),
    .out(\clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[10] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_fd_sc_hd__mux2_1 \clkgen.delay_155ns_2.genblk1[4].dly_binary.out_mux  (.A0(\clkgen.delay_155ns_2.genblk1[4].dly_binary.signal_w[16] ),
    .A1(\clkgen.delay_155ns_2.genblk1[3].dly_binary.out ),
    .S(\clkgen.delay_155ns_2.genblk1[4].dly_binary.bypass_in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.clk_dig_delayed_w ));
 sky130_fd_sc_hd__buf_4 \clkgen.delay_155ns_3.enablebuffer  (.A(enable_dlycontrol_in),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_3.enable_dlycontrol_w ));
 sky130_fd_sc_hd__and2_1 \clkgen.delay_155ns_3.genblk1[0].bypass_enable  (.A(\clkgen.delay_155ns_3.enable_dlycontrol_w ),
    .B(\clkgen.delay_155ns_3.bypass_enable_w[0] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_3.genblk1[0].dly_binary.bypass_in ));
 sky130_fd_sc_hd__inv_2 \clkgen.delay_155ns_3.genblk1[0].control_invert  (.A(dlycontrol3_in[0]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(\clkgen.delay_155ns_3.bypass_enable_w[0] ));
 sky130_fd_sc_hd__and2b_1 \clkgen.delay_155ns_3.genblk1[0].dly_binary.and_bypass_switch  (.A_N(\clkgen.delay_155ns_3.genblk1[0].dly_binary.bypass_in ),
    .B(\clkgen.delay_155ns_3.genblk1[0].dly_binary.in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_3.genblk1[0].dly_binary.signal_w[0] ));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_3.genblk1[0].dly_binary.genblk1[0].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_3.genblk1[0].dly_binary.signal_w[0] ),
    .out(\clkgen.delay_155ns_3.genblk1[0].dly_binary.signal_w[1] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_fd_sc_hd__mux2_1 \clkgen.delay_155ns_3.genblk1[0].dly_binary.out_mux  (.A0(\clkgen.delay_155ns_3.genblk1[0].dly_binary.signal_w[1] ),
    .A1(\clkgen.delay_155ns_3.genblk1[0].dly_binary.in ),
    .S(\clkgen.delay_155ns_3.genblk1[0].dly_binary.bypass_in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_3.genblk1[0].dly_binary.out ));
 sky130_fd_sc_hd__and2_1 \clkgen.delay_155ns_3.genblk1[1].bypass_enable  (.A(\clkgen.delay_155ns_3.enable_dlycontrol_w ),
    .B(\clkgen.delay_155ns_3.bypass_enable_w[1] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_3.genblk1[1].dly_binary.bypass_in ));
 sky130_fd_sc_hd__inv_2 \clkgen.delay_155ns_3.genblk1[1].control_invert  (.A(dlycontrol3_in[1]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(\clkgen.delay_155ns_3.bypass_enable_w[1] ));
 sky130_fd_sc_hd__and2b_1 \clkgen.delay_155ns_3.genblk1[1].dly_binary.and_bypass_switch  (.A_N(\clkgen.delay_155ns_3.genblk1[1].dly_binary.bypass_in ),
    .B(\clkgen.delay_155ns_3.genblk1[0].dly_binary.out ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_3.genblk1[1].dly_binary.signal_w[0] ));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_3.genblk1[1].dly_binary.genblk1[0].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_3.genblk1[1].dly_binary.signal_w[0] ),
    .out(\clkgen.delay_155ns_3.genblk1[1].dly_binary.signal_w[1] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_3.genblk1[1].dly_binary.genblk1[1].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_3.genblk1[1].dly_binary.signal_w[1] ),
    .out(\clkgen.delay_155ns_3.genblk1[1].dly_binary.signal_w[2] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_fd_sc_hd__mux2_1 \clkgen.delay_155ns_3.genblk1[1].dly_binary.out_mux  (.A0(\clkgen.delay_155ns_3.genblk1[1].dly_binary.signal_w[2] ),
    .A1(\clkgen.delay_155ns_3.genblk1[0].dly_binary.out ),
    .S(\clkgen.delay_155ns_3.genblk1[1].dly_binary.bypass_in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_3.genblk1[1].dly_binary.out ));
 sky130_fd_sc_hd__and2_1 \clkgen.delay_155ns_3.genblk1[2].bypass_enable  (.A(\clkgen.delay_155ns_3.enable_dlycontrol_w ),
    .B(\clkgen.delay_155ns_3.bypass_enable_w[2] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_3.genblk1[2].dly_binary.bypass_in ));
 sky130_fd_sc_hd__inv_2 \clkgen.delay_155ns_3.genblk1[2].control_invert  (.A(dlycontrol3_in[2]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(\clkgen.delay_155ns_3.bypass_enable_w[2] ));
 sky130_fd_sc_hd__and2b_1 \clkgen.delay_155ns_3.genblk1[2].dly_binary.and_bypass_switch  (.A_N(\clkgen.delay_155ns_3.genblk1[2].dly_binary.bypass_in ),
    .B(\clkgen.delay_155ns_3.genblk1[1].dly_binary.out ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_3.genblk1[2].dly_binary.signal_w[0] ));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_3.genblk1[2].dly_binary.genblk1[0].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_3.genblk1[2].dly_binary.signal_w[0] ),
    .out(\clkgen.delay_155ns_3.genblk1[2].dly_binary.signal_w[1] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_3.genblk1[2].dly_binary.genblk1[1].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_3.genblk1[2].dly_binary.signal_w[1] ),
    .out(\clkgen.delay_155ns_3.genblk1[2].dly_binary.signal_w[2] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_3.genblk1[2].dly_binary.genblk1[2].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_3.genblk1[2].dly_binary.signal_w[2] ),
    .out(\clkgen.delay_155ns_3.genblk1[2].dly_binary.signal_w[3] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_3.genblk1[2].dly_binary.genblk1[3].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_3.genblk1[2].dly_binary.signal_w[3] ),
    .out(\clkgen.delay_155ns_3.genblk1[2].dly_binary.signal_w[4] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_fd_sc_hd__mux2_1 \clkgen.delay_155ns_3.genblk1[2].dly_binary.out_mux  (.A0(\clkgen.delay_155ns_3.genblk1[2].dly_binary.signal_w[4] ),
    .A1(\clkgen.delay_155ns_3.genblk1[1].dly_binary.out ),
    .S(\clkgen.delay_155ns_3.genblk1[2].dly_binary.bypass_in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_3.genblk1[2].dly_binary.out ));
 sky130_fd_sc_hd__and2_1 \clkgen.delay_155ns_3.genblk1[3].bypass_enable  (.A(\clkgen.delay_155ns_3.enable_dlycontrol_w ),
    .B(\clkgen.delay_155ns_3.bypass_enable_w[3] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_3.genblk1[3].dly_binary.bypass_in ));
 sky130_fd_sc_hd__inv_2 \clkgen.delay_155ns_3.genblk1[3].control_invert  (.A(dlycontrol3_in[3]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(\clkgen.delay_155ns_3.bypass_enable_w[3] ));
 sky130_fd_sc_hd__and2b_1 \clkgen.delay_155ns_3.genblk1[3].dly_binary.and_bypass_switch  (.A_N(\clkgen.delay_155ns_3.genblk1[3].dly_binary.bypass_in ),
    .B(\clkgen.delay_155ns_3.genblk1[2].dly_binary.out ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_3.genblk1[3].dly_binary.signal_w[0] ));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_3.genblk1[3].dly_binary.genblk1[0].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_3.genblk1[3].dly_binary.signal_w[0] ),
    .out(\clkgen.delay_155ns_3.genblk1[3].dly_binary.signal_w[1] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_3.genblk1[3].dly_binary.genblk1[1].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_3.genblk1[3].dly_binary.signal_w[1] ),
    .out(\clkgen.delay_155ns_3.genblk1[3].dly_binary.signal_w[2] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_3.genblk1[3].dly_binary.genblk1[2].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_3.genblk1[3].dly_binary.signal_w[2] ),
    .out(\clkgen.delay_155ns_3.genblk1[3].dly_binary.signal_w[3] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_3.genblk1[3].dly_binary.genblk1[3].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_3.genblk1[3].dly_binary.signal_w[3] ),
    .out(\clkgen.delay_155ns_3.genblk1[3].dly_binary.signal_w[4] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_3.genblk1[3].dly_binary.genblk1[4].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_3.genblk1[3].dly_binary.signal_w[4] ),
    .out(\clkgen.delay_155ns_3.genblk1[3].dly_binary.signal_w[5] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_3.genblk1[3].dly_binary.genblk1[5].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_3.genblk1[3].dly_binary.signal_w[5] ),
    .out(\clkgen.delay_155ns_3.genblk1[3].dly_binary.signal_w[6] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_3.genblk1[3].dly_binary.genblk1[6].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_3.genblk1[3].dly_binary.signal_w[6] ),
    .out(\clkgen.delay_155ns_3.genblk1[3].dly_binary.signal_w[7] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_3.genblk1[3].dly_binary.genblk1[7].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_3.genblk1[3].dly_binary.signal_w[7] ),
    .out(\clkgen.delay_155ns_3.genblk1[3].dly_binary.signal_w[8] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_fd_sc_hd__mux2_1 \clkgen.delay_155ns_3.genblk1[3].dly_binary.out_mux  (.A0(\clkgen.delay_155ns_3.genblk1[3].dly_binary.signal_w[8] ),
    .A1(\clkgen.delay_155ns_3.genblk1[2].dly_binary.out ),
    .S(\clkgen.delay_155ns_3.genblk1[3].dly_binary.bypass_in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_3.genblk1[3].dly_binary.out ));
 sky130_fd_sc_hd__and2_1 \clkgen.delay_155ns_3.genblk1[4].bypass_enable  (.A(\clkgen.delay_155ns_3.enable_dlycontrol_w ),
    .B(\clkgen.delay_155ns_3.bypass_enable_w[4] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_3.genblk1[4].dly_binary.bypass_in ));
 sky130_fd_sc_hd__inv_2 \clkgen.delay_155ns_3.genblk1[4].control_invert  (.A(dlycontrol3_in[4]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(\clkgen.delay_155ns_3.bypass_enable_w[4] ));
 sky130_fd_sc_hd__and2b_1 \clkgen.delay_155ns_3.genblk1[4].dly_binary.and_bypass_switch  (.A_N(\clkgen.delay_155ns_3.genblk1[4].dly_binary.bypass_in ),
    .B(\clkgen.delay_155ns_3.genblk1[3].dly_binary.out ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[0] ));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_3.genblk1[4].dly_binary.genblk1[0].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[0] ),
    .out(\clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[1] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_3.genblk1[4].dly_binary.genblk1[10].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[10] ),
    .out(\clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[11] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_3.genblk1[4].dly_binary.genblk1[11].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[11] ),
    .out(\clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[12] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_3.genblk1[4].dly_binary.genblk1[12].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[12] ),
    .out(\clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[13] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_3.genblk1[4].dly_binary.genblk1[13].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[13] ),
    .out(\clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[14] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_3.genblk1[4].dly_binary.genblk1[14].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[14] ),
    .out(\clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[15] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_3.genblk1[4].dly_binary.genblk1[15].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[15] ),
    .out(\clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[16] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_3.genblk1[4].dly_binary.genblk1[1].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[1] ),
    .out(\clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[2] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_3.genblk1[4].dly_binary.genblk1[2].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[2] ),
    .out(\clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[3] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_3.genblk1[4].dly_binary.genblk1[3].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[3] ),
    .out(\clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[4] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_3.genblk1[4].dly_binary.genblk1[4].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[4] ),
    .out(\clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[5] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_3.genblk1[4].dly_binary.genblk1[5].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[5] ),
    .out(\clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[6] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_3.genblk1[4].dly_binary.genblk1[6].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[6] ),
    .out(\clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[7] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_3.genblk1[4].dly_binary.genblk1[7].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[7] ),
    .out(\clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[8] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_3.genblk1[4].dly_binary.genblk1[8].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[8] ),
    .out(\clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[9] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \clkgen.delay_155ns_3.genblk1[4].dly_binary.genblk1[9].delay_unit  (.VPWR(VDD),
    .in(\clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[9] ),
    .out(\clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[10] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_fd_sc_hd__mux2_1 \clkgen.delay_155ns_3.genblk1[4].dly_binary.out_mux  (.A0(\clkgen.delay_155ns_3.genblk1[4].dly_binary.signal_w[16] ),
    .A1(\clkgen.delay_155ns_3.genblk1[3].dly_binary.out ),
    .S(\clkgen.delay_155ns_3.genblk1[4].dly_binary.bypass_in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.clk_comp_out ));
 sky130_fd_sc_hd__nor2b_1 \clkgen.nor1  (.A(\clkgen.clk_dig_delayed_w ),
    .B_N(\clkgen.enable_loop_in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(\clkgen.delay_155ns_3.genblk1[0].dly_binary.in ));
 sky130_mm_sc_hd_dlyPoly5ns delay_sample_n12 (.VPWR(VDD),
    .in(sample_n_in),
    .out(sample_n_1),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns delay_sample_p11 (.VPWR(VDD),
    .in(sample_p_in),
    .out(sample_p_1),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_fd_sc_hd__buf_4 \edgedetect.dly_315ns_1.enablebuffer  (.A(enable_dlycontrol_in),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\edgedetect.dly_315ns_1.enable_dlycontrol_w ));
 sky130_fd_sc_hd__and2_1 \edgedetect.dly_315ns_1.genblk1[0].bypass_enable  (.A(\edgedetect.dly_315ns_1.enable_dlycontrol_w ),
    .B(\edgedetect.dly_315ns_1.bypass_enable_w[0] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\edgedetect.dly_315ns_1.genblk1[0].dly_binary.bypass_in ));
 sky130_fd_sc_hd__inv_2 \edgedetect.dly_315ns_1.genblk1[0].control_invert  (.A(dlycontrol4_in[0]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(\edgedetect.dly_315ns_1.bypass_enable_w[0] ));
 sky130_fd_sc_hd__and2b_1 \edgedetect.dly_315ns_1.genblk1[0].dly_binary.and_bypass_switch  (.A_N(\edgedetect.dly_315ns_1.genblk1[0].dly_binary.bypass_in ),
    .B(\edgedetect.dly_315ns_1.genblk1[0].dly_binary.in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\edgedetect.dly_315ns_1.genblk1[0].dly_binary.signal_w[0] ));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[0].dly_binary.genblk1[0].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[0].dly_binary.signal_w[0] ),
    .out(\edgedetect.dly_315ns_1.genblk1[0].dly_binary.signal_w[1] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_fd_sc_hd__mux2_1 \edgedetect.dly_315ns_1.genblk1[0].dly_binary.out_mux  (.A0(\edgedetect.dly_315ns_1.genblk1[0].dly_binary.signal_w[1] ),
    .A1(\edgedetect.dly_315ns_1.genblk1[0].dly_binary.in ),
    .S(\edgedetect.dly_315ns_1.genblk1[0].dly_binary.bypass_in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\edgedetect.dly_315ns_1.genblk1[0].dly_binary.out ));
 sky130_fd_sc_hd__and2_1 \edgedetect.dly_315ns_1.genblk1[1].bypass_enable  (.A(\edgedetect.dly_315ns_1.enable_dlycontrol_w ),
    .B(\edgedetect.dly_315ns_1.bypass_enable_w[1] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\edgedetect.dly_315ns_1.genblk1[1].dly_binary.bypass_in ));
 sky130_fd_sc_hd__inv_2 \edgedetect.dly_315ns_1.genblk1[1].control_invert  (.A(dlycontrol4_in[1]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(\edgedetect.dly_315ns_1.bypass_enable_w[1] ));
 sky130_fd_sc_hd__and2b_1 \edgedetect.dly_315ns_1.genblk1[1].dly_binary.and_bypass_switch  (.A_N(\edgedetect.dly_315ns_1.genblk1[1].dly_binary.bypass_in ),
    .B(\edgedetect.dly_315ns_1.genblk1[0].dly_binary.out ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\edgedetect.dly_315ns_1.genblk1[1].dly_binary.signal_w[0] ));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[1].dly_binary.genblk1[0].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[1].dly_binary.signal_w[0] ),
    .out(\edgedetect.dly_315ns_1.genblk1[1].dly_binary.signal_w[1] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[1].dly_binary.genblk1[1].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[1].dly_binary.signal_w[1] ),
    .out(\edgedetect.dly_315ns_1.genblk1[1].dly_binary.signal_w[2] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_fd_sc_hd__mux2_1 \edgedetect.dly_315ns_1.genblk1[1].dly_binary.out_mux  (.A0(\edgedetect.dly_315ns_1.genblk1[1].dly_binary.signal_w[2] ),
    .A1(\edgedetect.dly_315ns_1.genblk1[0].dly_binary.out ),
    .S(\edgedetect.dly_315ns_1.genblk1[1].dly_binary.bypass_in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\edgedetect.dly_315ns_1.genblk1[1].dly_binary.out ));
 sky130_fd_sc_hd__and2_1 \edgedetect.dly_315ns_1.genblk1[2].bypass_enable  (.A(\edgedetect.dly_315ns_1.enable_dlycontrol_w ),
    .B(\edgedetect.dly_315ns_1.bypass_enable_w[2] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\edgedetect.dly_315ns_1.genblk1[2].dly_binary.bypass_in ));
 sky130_fd_sc_hd__inv_2 \edgedetect.dly_315ns_1.genblk1[2].control_invert  (.A(dlycontrol4_in[2]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(\edgedetect.dly_315ns_1.bypass_enable_w[2] ));
 sky130_fd_sc_hd__and2b_1 \edgedetect.dly_315ns_1.genblk1[2].dly_binary.and_bypass_switch  (.A_N(\edgedetect.dly_315ns_1.genblk1[2].dly_binary.bypass_in ),
    .B(\edgedetect.dly_315ns_1.genblk1[1].dly_binary.out ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\edgedetect.dly_315ns_1.genblk1[2].dly_binary.signal_w[0] ));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[2].dly_binary.genblk1[0].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[2].dly_binary.signal_w[0] ),
    .out(\edgedetect.dly_315ns_1.genblk1[2].dly_binary.signal_w[1] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[2].dly_binary.genblk1[1].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[2].dly_binary.signal_w[1] ),
    .out(\edgedetect.dly_315ns_1.genblk1[2].dly_binary.signal_w[2] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[2].dly_binary.genblk1[2].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[2].dly_binary.signal_w[2] ),
    .out(\edgedetect.dly_315ns_1.genblk1[2].dly_binary.signal_w[3] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[2].dly_binary.genblk1[3].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[2].dly_binary.signal_w[3] ),
    .out(\edgedetect.dly_315ns_1.genblk1[2].dly_binary.signal_w[4] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_fd_sc_hd__mux2_1 \edgedetect.dly_315ns_1.genblk1[2].dly_binary.out_mux  (.A0(\edgedetect.dly_315ns_1.genblk1[2].dly_binary.signal_w[4] ),
    .A1(\edgedetect.dly_315ns_1.genblk1[1].dly_binary.out ),
    .S(\edgedetect.dly_315ns_1.genblk1[2].dly_binary.bypass_in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\edgedetect.dly_315ns_1.genblk1[2].dly_binary.out ));
 sky130_fd_sc_hd__and2_1 \edgedetect.dly_315ns_1.genblk1[3].bypass_enable  (.A(\edgedetect.dly_315ns_1.enable_dlycontrol_w ),
    .B(\edgedetect.dly_315ns_1.bypass_enable_w[3] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\edgedetect.dly_315ns_1.genblk1[3].dly_binary.bypass_in ));
 sky130_fd_sc_hd__inv_2 \edgedetect.dly_315ns_1.genblk1[3].control_invert  (.A(dlycontrol4_in[3]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(\edgedetect.dly_315ns_1.bypass_enable_w[3] ));
 sky130_fd_sc_hd__and2b_1 \edgedetect.dly_315ns_1.genblk1[3].dly_binary.and_bypass_switch  (.A_N(\edgedetect.dly_315ns_1.genblk1[3].dly_binary.bypass_in ),
    .B(\edgedetect.dly_315ns_1.genblk1[2].dly_binary.out ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\edgedetect.dly_315ns_1.genblk1[3].dly_binary.signal_w[0] ));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[3].dly_binary.genblk1[0].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[3].dly_binary.signal_w[0] ),
    .out(\edgedetect.dly_315ns_1.genblk1[3].dly_binary.signal_w[1] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[3].dly_binary.genblk1[1].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[3].dly_binary.signal_w[1] ),
    .out(\edgedetect.dly_315ns_1.genblk1[3].dly_binary.signal_w[2] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[3].dly_binary.genblk1[2].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[3].dly_binary.signal_w[2] ),
    .out(\edgedetect.dly_315ns_1.genblk1[3].dly_binary.signal_w[3] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[3].dly_binary.genblk1[3].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[3].dly_binary.signal_w[3] ),
    .out(\edgedetect.dly_315ns_1.genblk1[3].dly_binary.signal_w[4] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[3].dly_binary.genblk1[4].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[3].dly_binary.signal_w[4] ),
    .out(\edgedetect.dly_315ns_1.genblk1[3].dly_binary.signal_w[5] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[3].dly_binary.genblk1[5].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[3].dly_binary.signal_w[5] ),
    .out(\edgedetect.dly_315ns_1.genblk1[3].dly_binary.signal_w[6] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[3].dly_binary.genblk1[6].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[3].dly_binary.signal_w[6] ),
    .out(\edgedetect.dly_315ns_1.genblk1[3].dly_binary.signal_w[7] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[3].dly_binary.genblk1[7].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[3].dly_binary.signal_w[7] ),
    .out(\edgedetect.dly_315ns_1.genblk1[3].dly_binary.signal_w[8] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_fd_sc_hd__mux2_1 \edgedetect.dly_315ns_1.genblk1[3].dly_binary.out_mux  (.A0(\edgedetect.dly_315ns_1.genblk1[3].dly_binary.signal_w[8] ),
    .A1(\edgedetect.dly_315ns_1.genblk1[2].dly_binary.out ),
    .S(\edgedetect.dly_315ns_1.genblk1[3].dly_binary.bypass_in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\edgedetect.dly_315ns_1.genblk1[3].dly_binary.out ));
 sky130_fd_sc_hd__and2_1 \edgedetect.dly_315ns_1.genblk1[4].bypass_enable  (.A(\edgedetect.dly_315ns_1.enable_dlycontrol_w ),
    .B(\edgedetect.dly_315ns_1.bypass_enable_w[4] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\edgedetect.dly_315ns_1.genblk1[4].dly_binary.bypass_in ));
 sky130_fd_sc_hd__inv_2 \edgedetect.dly_315ns_1.genblk1[4].control_invert  (.A(dlycontrol4_in[4]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(\edgedetect.dly_315ns_1.bypass_enable_w[4] ));
 sky130_fd_sc_hd__and2b_1 \edgedetect.dly_315ns_1.genblk1[4].dly_binary.and_bypass_switch  (.A_N(\edgedetect.dly_315ns_1.genblk1[4].dly_binary.bypass_in ),
    .B(\edgedetect.dly_315ns_1.genblk1[3].dly_binary.out ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[0] ));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[4].dly_binary.genblk1[0].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[0] ),
    .out(\edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[1] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[4].dly_binary.genblk1[10].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[10] ),
    .out(\edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[11] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[4].dly_binary.genblk1[11].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[11] ),
    .out(\edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[12] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[4].dly_binary.genblk1[12].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[12] ),
    .out(\edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[13] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[4].dly_binary.genblk1[13].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[13] ),
    .out(\edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[14] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[4].dly_binary.genblk1[14].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[14] ),
    .out(\edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[15] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[4].dly_binary.genblk1[15].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[15] ),
    .out(\edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[16] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[4].dly_binary.genblk1[1].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[1] ),
    .out(\edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[2] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[4].dly_binary.genblk1[2].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[2] ),
    .out(\edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[3] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[4].dly_binary.genblk1[3].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[3] ),
    .out(\edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[4] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[4].dly_binary.genblk1[4].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[4] ),
    .out(\edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[5] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[4].dly_binary.genblk1[5].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[5] ),
    .out(\edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[6] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[4].dly_binary.genblk1[6].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[6] ),
    .out(\edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[7] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[4].dly_binary.genblk1[7].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[7] ),
    .out(\edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[8] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[4].dly_binary.genblk1[8].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[8] ),
    .out(\edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[9] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[4].dly_binary.genblk1[9].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[9] ),
    .out(\edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[10] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_fd_sc_hd__mux2_1 \edgedetect.dly_315ns_1.genblk1[4].dly_binary.out_mux  (.A0(\edgedetect.dly_315ns_1.genblk1[4].dly_binary.signal_w[16] ),
    .A1(\edgedetect.dly_315ns_1.genblk1[3].dly_binary.out ),
    .S(\edgedetect.dly_315ns_1.genblk1[4].dly_binary.bypass_in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\edgedetect.dly_315ns_1.genblk1[4].dly_binary.out ));
 sky130_fd_sc_hd__and2_1 \edgedetect.dly_315ns_1.genblk1[5].bypass_enable  (.A(\edgedetect.dly_315ns_1.enable_dlycontrol_w ),
    .B(\edgedetect.dly_315ns_1.bypass_enable_w[5] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.bypass_in ));
 sky130_fd_sc_hd__inv_2 \edgedetect.dly_315ns_1.genblk1[5].control_invert  (.A(dlycontrol4_in[5]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(\edgedetect.dly_315ns_1.bypass_enable_w[5] ));
 sky130_fd_sc_hd__and2b_1 \edgedetect.dly_315ns_1.genblk1[5].dly_binary.and_bypass_switch  (.A_N(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.bypass_in ),
    .B(\edgedetect.dly_315ns_1.genblk1[4].dly_binary.out ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[0] ));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[5].dly_binary.genblk1[0].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[0] ),
    .out(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[1] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[5].dly_binary.genblk1[10].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[10] ),
    .out(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[11] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[5].dly_binary.genblk1[11].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[11] ),
    .out(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[12] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[5].dly_binary.genblk1[12].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[12] ),
    .out(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[13] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[5].dly_binary.genblk1[13].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[13] ),
    .out(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[14] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[5].dly_binary.genblk1[14].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[14] ),
    .out(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[15] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[5].dly_binary.genblk1[15].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[15] ),
    .out(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[16] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[5].dly_binary.genblk1[16].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[16] ),
    .out(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[17] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[5].dly_binary.genblk1[17].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[17] ),
    .out(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[18] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[5].dly_binary.genblk1[18].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[18] ),
    .out(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[19] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[5].dly_binary.genblk1[19].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[19] ),
    .out(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[20] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[5].dly_binary.genblk1[1].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[1] ),
    .out(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[2] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[5].dly_binary.genblk1[20].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[20] ),
    .out(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[21] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[5].dly_binary.genblk1[21].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[21] ),
    .out(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[22] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[5].dly_binary.genblk1[22].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[22] ),
    .out(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[23] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[5].dly_binary.genblk1[23].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[23] ),
    .out(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[24] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[5].dly_binary.genblk1[24].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[24] ),
    .out(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[25] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[5].dly_binary.genblk1[25].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[25] ),
    .out(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[26] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[5].dly_binary.genblk1[26].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[26] ),
    .out(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[27] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[5].dly_binary.genblk1[27].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[27] ),
    .out(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[28] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[5].dly_binary.genblk1[28].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[28] ),
    .out(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[29] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[5].dly_binary.genblk1[29].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[29] ),
    .out(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[30] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[5].dly_binary.genblk1[2].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[2] ),
    .out(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[3] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[5].dly_binary.genblk1[30].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[30] ),
    .out(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[31] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[5].dly_binary.genblk1[31].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[31] ),
    .out(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[32] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[5].dly_binary.genblk1[3].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[3] ),
    .out(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[4] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[5].dly_binary.genblk1[4].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[4] ),
    .out(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[5] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[5].dly_binary.genblk1[5].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[5] ),
    .out(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[6] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[5].dly_binary.genblk1[6].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[6] ),
    .out(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[7] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[5].dly_binary.genblk1[7].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[7] ),
    .out(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[8] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[5].dly_binary.genblk1[8].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[8] ),
    .out(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[9] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_mm_sc_hd_dlyPoly5ns \edgedetect.dly_315ns_1.genblk1[5].dly_binary.genblk1[9].delay_unit  (.VPWR(VDD),
    .in(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[9] ),
    .out(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[10] ),
    .VGND(VSS),
    .VPB(VDD),
    .VNB(VSS));
 sky130_fd_sc_hd__mux2_1 \edgedetect.dly_315ns_1.genblk1[5].dly_binary.out_mux  (.A0(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.signal_w[32] ),
    .A1(\edgedetect.dly_315ns_1.genblk1[4].dly_binary.out ),
    .S(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.bypass_in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.out ));
 sky130_fd_sc_hd__nor2b_1 \edgedetect.nor1  (.A(\edgedetect.dly_315ns_1.genblk1[5].dly_binary.out ),
    .B_N(\edgedetect.dly_315ns_1.genblk1[0].dly_binary.in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .Y(\edgedetect.start_conv_edge_w ));
 sky130_fd_sc_hd__or2_1 \edgedetect.or1  (.A(\edgedetect.start_conv_edge_w ),
    .B(\edgedetect.ena_in ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.enable_loop_in ));
 sky130_fd_sc_hd__buf_1 inbuf_1 (.A(ena_in),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\edgedetect.ena_in ));
 sky130_fd_sc_hd__buf_1 inbuf_2 (.A(start_conv_in),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\edgedetect.dly_315ns_1.genblk1[0].dly_binary.in ));
 sky130_fd_sc_hd__buf_1 inbuf_3 (.A(ndecision_finish_in),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(\clkgen.delay_155ns_1.genblk1[0].dly_binary.in ));
 sky130_fd_sc_hd__bufbuf_8 outbuf_1 (.A(\clkgen.clk_dig_out ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(clk_dig_out));
 sky130_fd_sc_hd__bufbuf_8 outbuf_2 (.A(\clkgen.clk_comp_out ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(clk_comp_out));
 sky130_fd_sc_hd__bufbuf_8 outbuf_3 (.A(sample_p_1),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(sample_p_out));
 sky130_fd_sc_hd__bufbuf_8 outbuf_4 (.A(sample_n_1),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VDD),
    .VPWR(VDD),
    .X(sample_n_out));
endmodule
